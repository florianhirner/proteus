`timescale 1ns / 1ps

//-------------------------------------------------------------------------------------------------

module tw_rom_0_ntt_nwc
#(
    parameter LOGN  = 0,
    parameter LOGQ  = 64,
    parameter DELAY = 1,
    parameter STAGE = 0
)(
    input            clk,
    input [LOGN-1:0] raddr,
    output[LOGQ-1:0] b
);

(* rom_style = "distributed" *)
reg [LOGQ-1:0] brom_out, brom_out2;

always @(posedge clk) begin
    case(raddr[0:0])
    1'd0: brom_out <= 64'd6551015095526749063;
    default: brom_out <= 64'h1;
    endcase
end

generate
    if(DELAY == 1) begin
        assign b = brom_out;
    end
endgenerate

endmodule

//-------------------------------------------------------------------------------------------------

module tw_rom_1_ntt_nwc
#(
    parameter LOGN  = 1,
    parameter LOGQ  = 64,
    parameter DELAY = 1,
    parameter STAGE = 1
)(
    input            clk,
    input [LOGN-1:0] raddr,
    output[LOGQ-1:0] b
);

(* rom_style = "distributed" *)
reg [LOGQ-1:0] brom_out, brom_out2;

always @(posedge clk) begin
    case(raddr[STAGE-1:0])
    2'd0: brom_out <= 64'd5976068779477487504;
    2'd1: brom_out <= 64'd3392617565049336557;
    default: brom_out <= 64'h1;
    endcase
end

generate
    if(DELAY == 1) begin
        assign b = brom_out;
    end
endgenerate

endmodule

//-------------------------------------------------------------------------------------------------

module tw_rom_2_ntt_nwc
#(
    parameter LOGN  = 2,
    parameter LOGQ  = 64,
    parameter DELAY = 1,
    parameter STAGE = 2
)(
    input            clk,
    input [LOGN-1:0] raddr,
    output[LOGQ-1:0] b
);

(* rom_style = "distributed" *)
reg [LOGQ-1:0] brom_out, brom_out2;

always @(posedge clk) begin
    case(raddr[STAGE-1:0])
    3'd0: brom_out <= 64'd2881966912403406253;
    3'd2: brom_out <= 64'd2991444385089030097;
    3'd1: brom_out <= 64'd5792979130194094298;
    3'd3: brom_out <= 64'd699101306064864663;
    default: brom_out <= 64'h1;
    endcase
end

generate
    if(DELAY == 1) begin
        assign b = brom_out;
    end
endgenerate

endmodule

//-------------------------------------------------------------------------------------------------

module tw_rom_3_ntt_nwc
#(
    parameter LOGN  = 3,
    parameter LOGQ  = 64,
    parameter DELAY = 1,
    parameter STAGE = 3
)(
    input            clk,
    input [LOGN-1:0] raddr,
    output[LOGQ-1:0] b
);

(* rom_style = "distributed" *)
reg [LOGQ-1:0] brom_out, brom_out2;

always @(posedge clk) begin
    case(raddr[STAGE-1:0])
    4'd0: brom_out <= 64'd5917339183240377480;
    4'd4: brom_out <= 64'd5908178380096272369;
    4'd2: brom_out <= 64'd4066724171054462909;
    4'd6: brom_out <= 64'd1002059954001900696;
    4'd1: brom_out <= 64'd7147821265559899415;
    4'd5: brom_out <= 64'd7646914504675205489;
    4'd3: brom_out <= 64'd2803267708398697040;
    4'd7: brom_out <= 64'd1670791095363685175;
    default: brom_out <= 64'h1;
    endcase
end

generate
    if(DELAY == 1) begin
        assign b = brom_out;
    end
endgenerate

endmodule

//-------------------------------------------------------------------------------------------------

module tw_rom_4_ntt_nwc
#(
    parameter LOGN  = 4,
    parameter LOGQ  = 64,
    parameter DELAY = 1,
    parameter STAGE = 4
)(
    input            clk,
    input [LOGN-1:0] raddr,
    output[LOGQ-1:0] b
);

(* rom_style = "distributed" *)
reg [LOGQ-1:0] brom_out, brom_out2;

always @(posedge clk) begin
    case(raddr[STAGE-1:0])
    5'd0: brom_out <= 64'd8706294438413809553;
    5'd8: brom_out <= 64'd8872444489401680815;
    5'd4: brom_out <= 64'd3874323780530106533;
    5'd12: brom_out <= 64'd5039744181953194803;
    5'd2: brom_out <= 64'd1624553938728686361;
    5'd10: brom_out <= 64'd9166670786663116443;
    5'd6: brom_out <= 64'd2737158020017696281;
    5'd14: brom_out <= 64'd7923677684682802987;
    5'd1: brom_out <= 64'd4110363107264655732;
    5'd9: brom_out <= 64'd3547627594494878621;
    5'd5: brom_out <= 64'd2637886143940526168;
    5'd13: brom_out <= 64'd9185509849420767578;
    5'd3: brom_out <= 64'd3044098306375364542;
    5'd11: brom_out <= 64'd4393262027419573708;
    5'd7: brom_out <= 64'd1065160304167154726;
    5'd15: brom_out <= 64'd228503451388919711;
    default: brom_out <= 64'h1;
    endcase
end

generate
    if(DELAY == 1) begin
        assign b = brom_out;
    end
endgenerate

endmodule

//-------------------------------------------------------------------------------------------------

module tw_rom_5_ntt_nwc
#(
    parameter LOGN  = 5,
    parameter LOGQ  = 64,
    parameter DELAY = 1,
    parameter STAGE = 5
)(
    input            clk,
    input [LOGN-1:0] raddr,
    output[LOGQ-1:0] b
);

(* rom_style = "distributed" *)
reg [LOGQ-1:0] brom_out, brom_out2;

always @(posedge clk) begin
    case(raddr[STAGE-1:0])
    6'd0: brom_out <= 64'd6984365454624050605;
    6'd16: brom_out <= 64'd284038871857826017;
    6'd8: brom_out <= 64'd8439932809411290039;
    6'd24: brom_out <= 64'd8216761589456164;
    6'd4: brom_out <= 64'd735439083491420630;
    6'd20: brom_out <= 64'd8124953238658307565;
    6'd12: brom_out <= 64'd5596038778869841895;
    6'd28: brom_out <= 64'd69843017785227084;
    6'd2: brom_out <= 64'd3950921523134993168;
    6'd18: brom_out <= 64'd1687335542159875606;
    6'd10: brom_out <= 64'd8309796333647791448;
    6'd26: brom_out <= 64'd4836003352449041316;
    6'd6: brom_out <= 64'd8826561644056073004;
    6'd22: brom_out <= 64'd2141707773911427712;
    6'd14: brom_out <= 64'd3003943219615574075;
    6'd30: brom_out <= 64'd8823464365455855293;
    6'd1: brom_out <= 64'd6158485483849164736;
    6'd17: brom_out <= 64'd2669547459691193432;
    6'd9: brom_out <= 64'd1085106348447748099;
    6'd25: brom_out <= 64'd1628906345678539120;
    6'd5: brom_out <= 64'd5875474638474206446;
    6'd21: brom_out <= 64'd5654726277541044038;
    6'd13: brom_out <= 64'd6071971305117248446;
    6'd29: brom_out <= 64'd5126845061066175356;
    6'd3: brom_out <= 64'd2194362728065833183;
    6'd19: brom_out <= 64'd2468663283803736374;
    6'd11: brom_out <= 64'd4291000205908552613;
    6'd27: brom_out <= 64'd9003279055065478956;
    6'd7: brom_out <= 64'd3522401398456133729;
    6'd23: brom_out <= 64'd5729951333194461427;
    6'd15: brom_out <= 64'd4910995540748981844;
    6'd31: brom_out <= 64'd700730835196570872;
    default: brom_out <= 64'h1;
    endcase
end

generate
    if(DELAY == 1) begin
        assign b = brom_out;
    end
endgenerate

endmodule

//-------------------------------------------------------------------------------------------------

module tw_rom_6_ntt_nwc
#(
    parameter LOGN  = 6,
    parameter LOGQ  = 64,
    parameter DELAY = 1,
    parameter STAGE = 6
)(
    input            clk,
    input [LOGN-1:0] raddr,
    output[LOGQ-1:0] b
);

(* rom_style = "distributed" *)
reg [LOGQ-1:0] brom_out, brom_out2;

always @(posedge clk) begin
    case(raddr[STAGE-1:0])
    7'd0: brom_out <= 64'd269998454485676360;
    7'd32: brom_out <= 64'd4040899244153570090;
    7'd16: brom_out <= 64'd1271675644934090509;
    7'd48: brom_out <= 64'd2263269548655216762;
    7'd8: brom_out <= 64'd1219064800028085468;
    7'd40: brom_out <= 64'd6281663284576107517;
    7'd24: brom_out <= 64'd5318975219191802577;
    7'd56: brom_out <= 64'd5893272571222366297;
    7'd4: brom_out <= 64'd8174323033676948403;
    7'd36: brom_out <= 64'd9076916340755116149;
    7'd20: brom_out <= 64'd4710964611444245301;
    7'd52: brom_out <= 64'd307156682351195017;
    7'd12: brom_out <= 64'd4717392765204693644;
    7'd44: brom_out <= 64'd1555308162728177297;
    7'd28: brom_out <= 64'd4083878445077305523;
    7'd60: brom_out <= 64'd3280526131456603436;
    7'd2: brom_out <= 64'd6626061600160634657;
    7'd34: brom_out <= 64'd2703826489472427745;
    7'd18: brom_out <= 64'd4363004334232094865;
    7'd50: brom_out <= 64'd5471972468712594632;
    7'd10: brom_out <= 64'd2926075365041679386;
    7'd42: brom_out <= 64'd3115848091286679823;
    7'd26: brom_out <= 64'd2216455649141208680;
    7'd58: brom_out <= 64'd375356035198548383;
    7'd6: brom_out <= 64'd8070303386396255336;
    7'd38: brom_out <= 64'd5944864576936445287;
    7'd22: brom_out <= 64'd7086452204833135780;
    7'd54: brom_out <= 64'd7995675456769788758;
    7'd14: brom_out <= 64'd221168427156668620;
    7'd46: brom_out <= 64'd4919595983980879989;
    7'd30: brom_out <= 64'd3598379093835291182;
    7'd62: brom_out <= 64'd7002130558985726630;
    7'd1: brom_out <= 64'd5653377166457707394;
    7'd33: brom_out <= 64'd2529239563039080875;
    7'd17: brom_out <= 64'd9036648888917473750;
    7'd49: brom_out <= 64'd8186964208105355814;
    7'd9: brom_out <= 64'd544940125055465581;
    7'd41: brom_out <= 64'd5782598045554155253;
    7'd25: brom_out <= 64'd6458351418566661432;
    7'd57: brom_out <= 64'd7645071031480098655;
    7'd5: brom_out <= 64'd4573453364429337213;
    7'd37: brom_out <= 64'd4938289008039594695;
    7'd21: brom_out <= 64'd4441590473776765300;
    7'd53: brom_out <= 64'd6436331060924184539;
    7'd13: brom_out <= 64'd3526492789053904424;
    7'd45: brom_out <= 64'd7010796944267998638;
    7'd29: brom_out <= 64'd6019869478886392755;
    7'd61: brom_out <= 64'd8323983203612776937;
    7'd3: brom_out <= 64'd7345482494331839697;
    7'd35: brom_out <= 64'd538390155169630246;
    7'd19: brom_out <= 64'd1403509903281381135;
    7'd51: brom_out <= 64'd3528090222809025860;
    7'd11: brom_out <= 64'd6222003843073247882;
    7'd43: brom_out <= 64'd3558399091024426444;
    7'd27: brom_out <= 64'd4050420130283138042;
    7'd59: brom_out <= 64'd796180145389681740;
    7'd7: brom_out <= 64'd6564530672913887453;
    7'd39: brom_out <= 64'd1178188298187125443;
    7'd23: brom_out <= 64'd6665838607271236324;
    7'd55: brom_out <= 64'd1827606411485443129;
    7'd15: brom_out <= 64'd9025502593406216690;
    7'd47: brom_out <= 64'd1376701315345052441;
    7'd31: brom_out <= 64'd8856063189815385885;
    7'd63: brom_out <= 64'd2113561489472542490;
    default: brom_out <= 64'h1;
    endcase
end

generate
    if(DELAY == 1) begin
        assign b = brom_out;
    end
endgenerate

endmodule

//-------------------------------------------------------------------------------------------------

module tw_rom_7_ntt_nwc
#(
    parameter LOGN  = 7,
    parameter LOGQ  = 64,
    parameter DELAY = 1,
    parameter STAGE = 7
)(
    input            clk,
    input [LOGN-1:0] raddr,
    output[LOGQ-1:0] b
);

(* rom_style = "distributed" *)
reg [LOGQ-1:0] brom_out, brom_out2;

always @(posedge clk) begin
    case(raddr[STAGE-1:0])
    8'd0: brom_out <= 64'd1299456045732977605;
    8'd64: brom_out <= 64'd3796382495133268725;
    8'd32: brom_out <= 64'd593042282816257658;
    8'd96: brom_out <= 64'd7479147464852913991;
    8'd16: brom_out <= 64'd8852621130615879035;
    8'd80: brom_out <= 64'd1122397655549924356;
    8'd48: brom_out <= 64'd222968537858942369;
    8'd112: brom_out <= 64'd8219959792660589692;
    8'd8: brom_out <= 64'd3561119328844693546;
    8'd72: brom_out <= 64'd4682857295746554344;
    8'd40: brom_out <= 64'd3603203538984367077;
    8'd104: brom_out <= 64'd1490887556607246244;
    8'd24: brom_out <= 64'd3149227341269420724;
    8'd88: brom_out <= 64'd3065938557921374089;
    8'd56: brom_out <= 64'd1618067356643750162;
    8'd120: brom_out <= 64'd5989914729659460893;
    8'd4: brom_out <= 64'd1984480336129885140;
    8'd68: brom_out <= 64'd4613289516563687559;
    8'd36: brom_out <= 64'd5718867093180509803;
    8'd100: brom_out <= 64'd3064309850488305304;
    8'd20: brom_out <= 64'd3586995478868233709;
    8'd84: brom_out <= 64'd7173654840489607776;
    8'd52: brom_out <= 64'd5607163649712091882;
    8'd116: brom_out <= 64'd2139689406997953411;
    8'd12: brom_out <= 64'd5233426006749936404;
    8'd76: brom_out <= 64'd57560180524151836;
    8'd44: brom_out <= 64'd5320908759602881481;
    8'd108: brom_out <= 64'd1546731779372361302;
    8'd28: brom_out <= 64'd7940586545958498989;
    8'd92: brom_out <= 64'd4159689793066360690;
    8'd60: brom_out <= 64'd8151167855892330172;
    8'd124: brom_out <= 64'd498968785704607628;
    8'd2: brom_out <= 64'd810060818546034655;
    8'd66: brom_out <= 64'd2554384204381077376;
    8'd34: brom_out <= 64'd9170359323010223211;
    8'd98: brom_out <= 64'd6925371594294004533;
    8'd18: brom_out <= 64'd4936662293846854616;
    8'd82: brom_out <= 64'd4625294087119433729;
    8'd50: brom_out <= 64'd3365288337767276247;
    8'd114: brom_out <= 64'd8225172405297280263;
    8'd10: brom_out <= 64'd3531419639158455240;
    8'd74: brom_out <= 64'd8818463071528412136;
    8'd42: brom_out <= 64'd5684075750352032262;
    8'd106: brom_out <= 64'd2923414615723271043;
    8'd26: brom_out <= 64'd7048641871031816;
    8'd90: brom_out <= 64'd5418439566171715291;
    8'd58: brom_out <= 64'd2803062370827609981;
    8'd122: brom_out <= 64'd5003529372930301250;
    8'd6: brom_out <= 64'd2808688244394002011;
    8'd70: brom_out <= 64'd8345571030034495946;
    8'd38: brom_out <= 64'd809486194630696952;
    8'd102: brom_out <= 64'd7705829573832500897;
    8'd22: brom_out <= 64'd7289325041362829578;
    8'd86: brom_out <= 64'd5208814341045079371;
    8'd54: brom_out <= 64'd2023644405886518221;
    8'd118: brom_out <= 64'd9162350688835803463;
    8'd14: brom_out <= 64'd240070673848085803;
    8'd78: brom_out <= 64'd1837680713908133646;
    8'd46: brom_out <= 64'd1232654478032123658;
    8'd110: brom_out <= 64'd869826359180825983;
    8'd30: brom_out <= 64'd7748187342122623094;
    8'd94: brom_out <= 64'd2240289491309476277;
    8'd62: brom_out <= 64'd9009408318896786413;
    8'd126: brom_out <= 64'd8584995141337045279;
    8'd1: brom_out <= 64'd9033387621081412018;
    8'd65: brom_out <= 64'd5683041679221725246;
    8'd33: brom_out <= 64'd1177438167634269823;
    8'd97: brom_out <= 64'd6982695801609760735;
    8'd17: brom_out <= 64'd1865389637899575391;
    8'd81: brom_out <= 64'd8697599446790123293;
    8'd49: brom_out <= 64'd5000944239179137954;
    8'd113: brom_out <= 64'd4439925312673350003;
    8'd9: brom_out <= 64'd2319035647868930894;
    8'd73: brom_out <= 64'd5040843640203270416;
    8'd41: brom_out <= 64'd6828380608571071779;
    8'd105: brom_out <= 64'd3107918471259441615;
    8'd25: brom_out <= 64'd4312120720500409507;
    8'd89: brom_out <= 64'd6550225160897858344;
    8'd57: brom_out <= 64'd7741923924364988008;
    8'd121: brom_out <= 64'd3615127351505505023;
    8'd5: brom_out <= 64'd6375267241083926885;
    8'd69: brom_out <= 64'd1952843272151728048;
    8'd37: brom_out <= 64'd7929071200947786101;
    8'd101: brom_out <= 64'd6626178562688381462;
    8'd21: brom_out <= 64'd5712154480457087476;
    8'd85: brom_out <= 64'd750361034814781007;
    8'd53: brom_out <= 64'd1455837426791755297;
    8'd117: brom_out <= 64'd511527761999251354;
    8'd13: brom_out <= 64'd5682374489572555945;
    8'd77: brom_out <= 64'd684639643803771175;
    8'd45: brom_out <= 64'd3372994486386929879;
    8'd109: brom_out <= 64'd4849682055056439114;
    8'd29: brom_out <= 64'd5446263128435942946;
    8'd93: brom_out <= 64'd4919750730687193807;
    8'd61: brom_out <= 64'd4667723862850537194;
    8'd125: brom_out <= 64'd7471415495952780188;
    8'd3: brom_out <= 64'd8914698016797979130;
    8'd67: brom_out <= 64'd9106909176665937792;
    8'd35: brom_out <= 64'd739218949392655402;
    8'd99: brom_out <= 64'd6849437044168275747;
    8'd19: brom_out <= 64'd1845447672304840611;
    8'd83: brom_out <= 64'd5991059833680697521;
    8'd51: brom_out <= 64'd5293457782313866956;
    8'd115: brom_out <= 64'd5173422508798334624;
    8'd11: brom_out <= 64'd3367056065757602806;
    8'd75: brom_out <= 64'd6574977840107373503;
    8'd43: brom_out <= 64'd6707938413484059878;
    8'd107: brom_out <= 64'd1641922973023157952;
    8'd27: brom_out <= 64'd5311697839062869272;
    8'd91: brom_out <= 64'd8692551628537520016;
    8'd59: brom_out <= 64'd5746142847633122703;
    8'd123: brom_out <= 64'd5423351720389833865;
    8'd7: brom_out <= 64'd8037037384829722617;
    8'd71: brom_out <= 64'd4078971191093288272;
    8'd39: brom_out <= 64'd4619323584991910886;
    8'd103: brom_out <= 64'd8798316185508471405;
    8'd23: brom_out <= 64'd616529505270125954;
    8'd87: brom_out <= 64'd4764036910647300995;
    8'd55: brom_out <= 64'd5243772136807645099;
    8'd119: brom_out <= 64'd4119508171639317112;
    8'd15: brom_out <= 64'd1907082839763808740;
    8'd79: brom_out <= 64'd5873106135293020355;
    8'd47: brom_out <= 64'd4070504440077246346;
    8'd111: brom_out <= 64'd7672998258368931866;
    8'd31: brom_out <= 64'd4533570374417505243;
    8'd95: brom_out <= 64'd5939667306004532036;
    8'd63: brom_out <= 64'd4891968351182874667;
    8'd127: brom_out <= 64'd7269045898348823146;
    default: brom_out <= 64'h1;
    endcase
end

generate
    if(DELAY == 1) begin
        assign b = brom_out;
    end
endgenerate

endmodule

//-------------------------------------------------------------------------------------------------

module tw_rom_8_ntt_nwc
#(
    parameter LOGN  = 8,
    parameter LOGQ  = 64,
    parameter DELAY = 1,
    parameter STAGE = 8
)(
    input            clk,
    input [LOGN-1:0] raddr,
    output[LOGQ-1:0] b
);

(* ram_style = "block" *)
reg [LOGQ-1:0] brom_out, brom_out2;

always @(posedge clk) begin
    case(raddr[STAGE-1:0])
    9'd0: brom_out <= 64'd7605493872853681221;
    9'd128: brom_out <= 64'd8652315721870189437;
    9'd64: brom_out <= 64'd6061870125418198147;
    9'd192: brom_out <= 64'd2230049327513614869;
    9'd32: brom_out <= 64'd2925409531261716840;
    9'd160: brom_out <= 64'd4183299227927339195;
    9'd96: brom_out <= 64'd4452291514428477137;
    9'd224: brom_out <= 64'd655123889431899961;
    9'd16: brom_out <= 64'd4392041727794040139;
    9'd144: brom_out <= 64'd7993813175591520204;
    9'd80: brom_out <= 64'd1611893969776626643;
    9'd208: brom_out <= 64'd2757773614559033666;
    9'd48: brom_out <= 64'd1598994064067110291;
    9'd176: brom_out <= 64'd5713577346046003020;
    9'd112: brom_out <= 64'd8376944661285632772;
    9'd240: brom_out <= 64'd6268445540391799960;
    9'd8: brom_out <= 64'd2509796222201502174;
    9'd136: brom_out <= 64'd2343344652186686753;
    9'd72: brom_out <= 64'd6928014622416298408;
    9'd200: brom_out <= 64'd3468732936118861906;
    9'd40: brom_out <= 64'd3012117742719754636;
    9'd168: brom_out <= 64'd7083423175763586691;
    9'd104: brom_out <= 64'd2487979883454043411;
    9'd232: brom_out <= 64'd2275953281661646751;
    9'd24: brom_out <= 64'd5549948750888088698;
    9'd152: brom_out <= 64'd1549287551893278911;
    9'd88: brom_out <= 64'd4132551802894357262;
    9'd216: brom_out <= 64'd6230952056441481807;
    9'd56: brom_out <= 64'd967392942188980461;
    9'd184: brom_out <= 64'd8893614490103508778;
    9'd120: brom_out <= 64'd6953881865491377297;
    9'd248: brom_out <= 64'd6913883903315781469;
    9'd4: brom_out <= 64'd2123066514724381883;
    9'd132: brom_out <= 64'd7096948766236504610;
    9'd68: brom_out <= 64'd8791519766434938211;
    9'd196: brom_out <= 64'd9102413699342598757;
    9'd36: brom_out <= 64'd5356334136853441455;
    9'd164: brom_out <= 64'd5808776274764837854;
    9'd100: brom_out <= 64'd7803653637595225642;
    9'd228: brom_out <= 64'd8247980103556855667;
    9'd20: brom_out <= 64'd2162992210110465427;
    9'd148: brom_out <= 64'd6854317339658753350;
    9'd84: brom_out <= 64'd7940540358792163042;
    9'd212: brom_out <= 64'd8051296741047110195;
    9'd52: brom_out <= 64'd6153283181782085767;
    9'd180: brom_out <= 64'd7593220218804307867;
    9'd116: brom_out <= 64'd1382872280811698552;
    9'd244: brom_out <= 64'd5139097896322553033;
    9'd12: brom_out <= 64'd1966154900029444318;
    9'd140: brom_out <= 64'd4585039786213636068;
    9'd76: brom_out <= 64'd853076967703601242;
    9'd204: brom_out <= 64'd4368700210148671551;
    9'd44: brom_out <= 64'd6548403254923287631;
    9'd172: brom_out <= 64'd4510264232516592952;
    9'd108: brom_out <= 64'd8108747189882628079;
    9'd236: brom_out <= 64'd6181066534637459237;
    9'd28: brom_out <= 64'd401958369407258982;
    9'd156: brom_out <= 64'd5798824876843371582;
    9'd92: brom_out <= 64'd7819977419197775899;
    9'd220: brom_out <= 64'd5011986474190685475;
    9'd60: brom_out <= 64'd6985849834050000541;
    9'd188: brom_out <= 64'd8743332571195579934;
    9'd124: brom_out <= 64'd6432548891759686389;
    9'd252: brom_out <= 64'd7087203385146507098;
    9'd2: brom_out <= 64'd7934371085285641861;
    9'd130: brom_out <= 64'd2240211916433264831;
    9'd66: brom_out <= 64'd8013822734360034103;
    9'd194: brom_out <= 64'd6798664954031634633;
    9'd34: brom_out <= 64'd543577740076728061;
    9'd162: brom_out <= 64'd7533491753178725717;
    9'd98: brom_out <= 64'd4110541742333500737;
    9'd226: brom_out <= 64'd2015889517693822068;
    9'd18: brom_out <= 64'd7153542761736184733;
    9'd146: brom_out <= 64'd5024898852976039286;
    9'd82: brom_out <= 64'd3118801396391702857;
    9'd210: brom_out <= 64'd8730278730941939396;
    9'd50: brom_out <= 64'd4359339040815035935;
    9'd178: brom_out <= 64'd220088159844794260;
    9'd114: brom_out <= 64'd6337223876791081151;
    9'd242: brom_out <= 64'd881381962624186811;
    9'd10: brom_out <= 64'd4332795524147639451;
    9'd138: brom_out <= 64'd3227682425404315158;
    9'd74: brom_out <= 64'd1021589499332145736;
    9'd202: brom_out <= 64'd8395167631823199941;
    9'd42: brom_out <= 64'd7993764406966422987;
    9'd170: brom_out <= 64'd5226535173943436928;
    9'd106: brom_out <= 64'd1314986123610772272;
    9'd234: brom_out <= 64'd4961919869715327681;
    9'd26: brom_out <= 64'd4346701462512900589;
    9'd154: brom_out <= 64'd5078991997579173257;
    9'd90: brom_out <= 64'd5695358218414993869;
    9'd218: brom_out <= 64'd198235807530720187;
    9'd58: brom_out <= 64'd6954602674252549157;
    9'd186: brom_out <= 64'd2816403948006974041;
    9'd122: brom_out <= 64'd3659981058207187100;
    9'd250: brom_out <= 64'd3016980039216328962;
    9'd6: brom_out <= 64'd2299841007653134372;
    9'd134: brom_out <= 64'd3847574256498121621;
    9'd70: brom_out <= 64'd994064848121607400;
    9'd198: brom_out <= 64'd1676869911627098617;
    9'd38: brom_out <= 64'd1297536695137410486;
    9'd166: brom_out <= 64'd7870108581299121483;
    9'd102: brom_out <= 64'd4456208975303951299;
    9'd230: brom_out <= 64'd5140288024937627165;
    9'd22: brom_out <= 64'd1287149587930120656;
    9'd150: brom_out <= 64'd3688954750038363726;
    9'd86: brom_out <= 64'd8634381596625442610;
    9'd214: brom_out <= 64'd6733707155866364304;
    9'd54: brom_out <= 64'd489108130890476637;
    9'd182: brom_out <= 64'd7135696680823117604;
    9'd118: brom_out <= 64'd6761610796267635122;
    9'd246: brom_out <= 64'd3740576396473059045;
    9'd14: brom_out <= 64'd299894953115934099;
    9'd142: brom_out <= 64'd1458993785378647509;
    9'd78: brom_out <= 64'd3510417462984237944;
    9'd206: brom_out <= 64'd1258669831230654444;
    9'd46: brom_out <= 64'd1990992240235617717;
    9'd174: brom_out <= 64'd1491544262489362891;
    9'd110: brom_out <= 64'd7977797132770592727;
    9'd238: brom_out <= 64'd6881112568257936145;
    9'd30: brom_out <= 64'd3098083654159802861;
    9'd158: brom_out <= 64'd3110559949174149380;
    9'd94: brom_out <= 64'd1297339388260599077;
    9'd222: brom_out <= 64'd6949147395764538964;
    9'd62: brom_out <= 64'd1744638522500329828;
    9'd190: brom_out <= 64'd3167756150689666531;
    9'd126: brom_out <= 64'd5590202575696230393;
    9'd254: brom_out <= 64'd3835383961103183096;
    9'd1: brom_out <= 64'd8213948439719346069;
    9'd129: brom_out <= 64'd15243861875148476;
    9'd65: brom_out <= 64'd5181330732459777477;
    9'd193: brom_out <= 64'd7538107808473199530;
    9'd33: brom_out <= 64'd270496797777326527;
    9'd161: brom_out <= 64'd2527297775950676908;
    9'd97: brom_out <= 64'd6650157038584548422;
    9'd225: brom_out <= 64'd8543830174923091154;
    9'd17: brom_out <= 64'd2908884142996516879;
    9'd145: brom_out <= 64'd8934879803166669689;
    9'd81: brom_out <= 64'd8041554051968754776;
    9'd209: brom_out <= 64'd7104811893195087792;
    9'd49: brom_out <= 64'd904660340594613265;
    9'd177: brom_out <= 64'd2744296939060575530;
    9'd113: brom_out <= 64'd2784388700362841711;
    9'd241: brom_out <= 64'd8498706274306490892;
    9'd9: brom_out <= 64'd7152306933764292478;
    9'd137: brom_out <= 64'd6832924728641330482;
    9'd73: brom_out <= 64'd8433488676012520446;
    9'd201: brom_out <= 64'd391518006782257654;
    9'd41: brom_out <= 64'd2057313745147478637;
    9'd169: brom_out <= 64'd1947243181919420491;
    9'd105: brom_out <= 64'd6229174968075775630;
    9'd233: brom_out <= 64'd3729764982569583119;
    9'd25: brom_out <= 64'd7125634071680409905;
    9'd153: brom_out <= 64'd7831437647304356508;
    9'd89: brom_out <= 64'd6222808144614635014;
    9'd217: brom_out <= 64'd1790792280522562723;
    9'd57: brom_out <= 64'd8888883322669091370;
    9'd185: brom_out <= 64'd654752926994167022;
    9'd121: brom_out <= 64'd4976637449741390052;
    9'd249: brom_out <= 64'd3083280881619226755;
    9'd5: brom_out <= 64'd8581206737579399620;
    9'd133: brom_out <= 64'd6463166748036722757;
    9'd69: brom_out <= 64'd4794628727443279888;
    9'd197: brom_out <= 64'd1568136098664689522;
    9'd37: brom_out <= 64'd5689831925774807956;
    9'd165: brom_out <= 64'd75966845172534173;
    9'd101: brom_out <= 64'd5892854050328892876;
    9'd229: brom_out <= 64'd976868090527140556;
    9'd21: brom_out <= 64'd6297866057014224030;
    9'd149: brom_out <= 64'd7284478466022368184;
    9'd85: brom_out <= 64'd6468256505106281226;
    9'd213: brom_out <= 64'd8026629062288902533;
    9'd53: brom_out <= 64'd3017602207931310620;
    9'd181: brom_out <= 64'd4249431574386262900;
    9'd117: brom_out <= 64'd7700372050315114363;
    9'd245: brom_out <= 64'd3363566323249637328;
    9'd13: brom_out <= 64'd7902540812321798218;
    9'd141: brom_out <= 64'd6017550373169230213;
    9'd77: brom_out <= 64'd6179534021270744021;
    9'd205: brom_out <= 64'd4934228471949137670;
    9'd45: brom_out <= 64'd1785088414017673288;
    9'd173: brom_out <= 64'd5551115908770807940;
    9'd109: brom_out <= 64'd6396414439770314375;
    9'd237: brom_out <= 64'd841949363898762459;
    9'd29: brom_out <= 64'd1427846036265206780;
    9'd157: brom_out <= 64'd2036591841189774695;
    9'd93: brom_out <= 64'd7099443897569798910;
    9'd221: brom_out <= 64'd6630229277550940928;
    9'd61: brom_out <= 64'd4187235956733982846;
    9'd189: brom_out <= 64'd2173356542276770935;
    9'd125: brom_out <= 64'd5184317378868141180;
    9'd253: brom_out <= 64'd6918964554399920495;
    9'd3: brom_out <= 64'd4765886196678305331;
    9'd131: brom_out <= 64'd8708624953667028585;
    9'd67: brom_out <= 64'd6903674494547403458;
    9'd195: brom_out <= 64'd6068442745462420874;
    9'd35: brom_out <= 64'd7923340214113792441;
    9'd163: brom_out <= 64'd235142833563334451;
    9'd99: brom_out <= 64'd1059548844895002697;
    9'd227: brom_out <= 64'd4798734633597747276;
    9'd19: brom_out <= 64'd5900439431409958858;
    9'd147: brom_out <= 64'd4506204908127599502;
    9'd83: brom_out <= 64'd8127637090793435339;
    9'd211: brom_out <= 64'd6460685242337216620;
    9'd51: brom_out <= 64'd749037117208255733;
    9'd179: brom_out <= 64'd5490294517849368108;
    9'd115: brom_out <= 64'd2215604315896092670;
    9'd243: brom_out <= 64'd6148609810148795929;
    9'd11: brom_out <= 64'd792297214988562254;
    9'd139: brom_out <= 64'd7104270022735541970;
    9'd75: brom_out <= 64'd2663302601066611311;
    9'd203: brom_out <= 64'd9209536114756024834;
    9'd43: brom_out <= 64'd3479065458090349436;
    9'd171: brom_out <= 64'd3592198641247208794;
    9'd107: brom_out <= 64'd1701272341948035267;
    9'd235: brom_out <= 64'd5412893724914022449;
    9'd27: brom_out <= 64'd173114810237193158;
    9'd155: brom_out <= 64'd3340259218302706899;
    9'd91: brom_out <= 64'd3022260544642597516;
    9'd219: brom_out <= 64'd9160052455972965925;
    9'd59: brom_out <= 64'd5301890443195662787;
    9'd187: brom_out <= 64'd4413826527383477878;
    9'd123: brom_out <= 64'd9119962653750090131;
    9'd251: brom_out <= 64'd9117660520541870682;
    9'd7: brom_out <= 64'd5779395201958353378;
    9'd135: brom_out <= 64'd111332146913263916;
    9'd71: brom_out <= 64'd7256022154194582960;
    9'd199: brom_out <= 64'd8444867741212273661;
    9'd39: brom_out <= 64'd2182902326656347159;
    9'd167: brom_out <= 64'd8100294372597586432;
    9'd103: brom_out <= 64'd2351375173829121150;
    9'd231: brom_out <= 64'd2600298912569494844;
    9'd23: brom_out <= 64'd3883460632785907410;
    9'd151: brom_out <= 64'd821107918729627811;
    9'd87: brom_out <= 64'd8077069361822515059;
    9'd215: brom_out <= 64'd4681773058202772675;
    9'd55: brom_out <= 64'd7009454947613216741;
    9'd183: brom_out <= 64'd4824069180043442917;
    9'd119: brom_out <= 64'd3130462232530454679;
    9'd247: brom_out <= 64'd5408302969401217960;
    9'd15: brom_out <= 64'd9104612624170912214;
    9'd143: brom_out <= 64'd4583234557640069978;
    9'd79: brom_out <= 64'd6415125647473131768;
    9'd207: brom_out <= 64'd6154077313509807261;
    9'd47: brom_out <= 64'd4535501105232824056;
    9'd175: brom_out <= 64'd9197868711120196895;
    9'd111: brom_out <= 64'd2314914454150418602;
    9'd239: brom_out <= 64'd4523573697502160143;
    9'd31: brom_out <= 64'd3031844387819961827;
    9'd159: brom_out <= 64'd8803778985884906727;
    9'd95: brom_out <= 64'd7603550242876584926;
    9'd223: brom_out <= 64'd7530731249570041776;
    9'd63: brom_out <= 64'd2914465977735506303;
    9'd191: brom_out <= 64'd2935114005611711057;
    9'd127: brom_out <= 64'd5145477708918912727;
    9'd255: brom_out <= 64'd8634110784643349010;
    default: brom_out <= 64'h1;
    endcase
end

generate
    if(DELAY == 1) begin
        assign b = brom_out;
    end
endgenerate

endmodule

//-------------------------------------------------------------------------------------------------

module tw_rom_9_ntt_nwc
#(
    parameter LOGN  = 9,
    parameter LOGQ  = 64,
    parameter DELAY = 1,
    parameter STAGE = 9
)(
    input            clk,
    input [LOGN-1:0] raddr,
    output[LOGQ-1:0] b
);

(* ram_style = "block" *)
reg [LOGQ-1:0] brom_out, brom_out2;

always @(posedge clk) begin
    case(raddr[STAGE-1:0])
    10'd0: brom_out <= 64'd6012871302989280084;
    10'd256: brom_out <= 64'd8288530531944855590;
    10'd128: brom_out <= 64'd6744020006969895307;
    10'd384: brom_out <= 64'd7131970059357333029;
    10'd64: brom_out <= 64'd9146187461299601623;
    10'd320: brom_out <= 64'd6427097281726706628;
    10'd192: brom_out <= 64'd1390063910113207289;
    10'd448: brom_out <= 64'd7889711590670918676;
    10'd32: brom_out <= 64'd8498480881154740865;
    10'd288: brom_out <= 64'd9103463721653978408;
    10'd160: brom_out <= 64'd548261701981485419;
    10'd416: brom_out <= 64'd4687421323741025393;
    10'd96: brom_out <= 64'd8249092968287330570;
    10'd352: brom_out <= 64'd8256294627998732981;
    10'd224: brom_out <= 64'd4568079005623157455;
    10'd480: brom_out <= 64'd3613147540994151386;
    10'd16: brom_out <= 64'd6756792246403704650;
    10'd272: brom_out <= 64'd6943865764417683064;
    10'd144: brom_out <= 64'd6351756831470743006;
    10'd400: brom_out <= 64'd637799399688374479;
    10'd80: brom_out <= 64'd2235543617824736075;
    10'd336: brom_out <= 64'd5395617652967469222;
    10'd208: brom_out <= 64'd6640287097552321424;
    10'd464: brom_out <= 64'd3815011943812575350;
    10'd48: brom_out <= 64'd4514892859148397044;
    10'd304: brom_out <= 64'd3136767173588347434;
    10'd176: brom_out <= 64'd7047875822701595031;
    10'd432: brom_out <= 64'd6282214430396223665;
    10'd112: brom_out <= 64'd3652792854953481228;
    10'd368: brom_out <= 64'd3058650903359729066;
    10'd240: brom_out <= 64'd8625960684678229166;
    10'd496: brom_out <= 64'd2939264214977633037;
    10'd8: brom_out <= 64'd2273617654662494576;
    10'd264: brom_out <= 64'd1445608483214028307;
    10'd136: brom_out <= 64'd5152644225124011089;
    10'd392: brom_out <= 64'd5266018003312504579;
    10'd72: brom_out <= 64'd8701208384429075876;
    10'd328: brom_out <= 64'd6514515671117556603;
    10'd200: brom_out <= 64'd1852954710699492504;
    10'd456: brom_out <= 64'd4891530948138436991;
    10'd40: brom_out <= 64'd2884516234218684811;
    10'd296: brom_out <= 64'd9135823465542849361;
    10'd168: brom_out <= 64'd6457789071063052555;
    10'd424: brom_out <= 64'd956565536080223686;
    10'd104: brom_out <= 64'd6492936536869808625;
    10'd360: brom_out <= 64'd635855831193566106;
    10'd232: brom_out <= 64'd47740789800497965;
    10'd488: brom_out <= 64'd5749262411298578370;
    10'd24: brom_out <= 64'd5266916899250488660;
    10'd280: brom_out <= 64'd1709606027938467824;
    10'd152: brom_out <= 64'd7280577718007746774;
    10'd408: brom_out <= 64'd1544674224130596118;
    10'd88: brom_out <= 64'd4515128673629883118;
    10'd344: brom_out <= 64'd5083175541303528685;
    10'd216: brom_out <= 64'd211205323560102598;
    10'd472: brom_out <= 64'd7984550382453767596;
    10'd56: brom_out <= 64'd7403262497201993765;
    10'd312: brom_out <= 64'd4585935009530136169;
    10'd184: brom_out <= 64'd7224435870105783327;
    10'd440: brom_out <= 64'd3820044292411662612;
    10'd120: brom_out <= 64'd4785516395754103712;
    10'd376: brom_out <= 64'd7978110531043641769;
    10'd248: brom_out <= 64'd3657039766247532725;
    10'd504: brom_out <= 64'd646297118098278772;
    10'd4: brom_out <= 64'd2564423744727517704;
    10'd260: brom_out <= 64'd4512365403662406081;
    10'd132: brom_out <= 64'd8522993162440537939;
    10'd388: brom_out <= 64'd3329822700088162495;
    10'd68: brom_out <= 64'd6306667576969932326;
    10'd324: brom_out <= 64'd4794722994419500598;
    10'd196: brom_out <= 64'd8995741913985100290;
    10'd452: brom_out <= 64'd7027244046667068898;
    10'd36: brom_out <= 64'd8346874721972884401;
    10'd292: brom_out <= 64'd6610810496821611972;
    10'd164: brom_out <= 64'd6926030477489072308;
    10'd420: brom_out <= 64'd4898893176619253892;
    10'd100: brom_out <= 64'd865268308687100412;
    10'd356: brom_out <= 64'd4054013996166535507;
    10'd228: brom_out <= 64'd2848313604941519881;
    10'd484: brom_out <= 64'd291195603844344417;
    10'd20: brom_out <= 64'd1408687539684857079;
    10'd276: brom_out <= 64'd3163609927867779470;
    10'd148: brom_out <= 64'd7137177962332868154;
    10'd404: brom_out <= 64'd8595678383967341286;
    10'd84: brom_out <= 64'd3516066647433260551;
    10'd340: brom_out <= 64'd8317588540207922448;
    10'd212: brom_out <= 64'd6796227057672368420;
    10'd468: brom_out <= 64'd1373369117410510866;
    10'd52: brom_out <= 64'd8117367890929318445;
    10'd308: brom_out <= 64'd978720527126678484;
    10'd180: brom_out <= 64'd1213734665504106333;
    10'd436: brom_out <= 64'd3111218648416961668;
    10'd116: brom_out <= 64'd7985210005529564458;
    10'd372: brom_out <= 64'd6301640391988730655;
    10'd244: brom_out <= 64'd3473787664538686576;
    10'd500: brom_out <= 64'd2804463966393397031;
    10'd12: brom_out <= 64'd2934009396408142147;
    10'd268: brom_out <= 64'd5407047594096528025;
    10'd140: brom_out <= 64'd8336322066205089657;
    10'd396: brom_out <= 64'd8817464271798224027;
    10'd76: brom_out <= 64'd2331992164875830888;
    10'd332: brom_out <= 64'd1141036854004408858;
    10'd204: brom_out <= 64'd2721341105491390085;
    10'd460: brom_out <= 64'd3868531777045828691;
    10'd44: brom_out <= 64'd6252329300465472480;
    10'd300: brom_out <= 64'd5802647509516054700;
    10'd172: brom_out <= 64'd787340924847783803;
    10'd428: brom_out <= 64'd5549270204663924183;
    10'd108: brom_out <= 64'd1097341705165972594;
    10'd364: brom_out <= 64'd3468411571066471426;
    10'd236: brom_out <= 64'd7140722186488696864;
    10'd492: brom_out <= 64'd2040235830658135393;
    10'd28: brom_out <= 64'd4218632253198916038;
    10'd284: brom_out <= 64'd7452519829483945138;
    10'd156: brom_out <= 64'd4551293125869120088;
    10'd412: brom_out <= 64'd1607600945152906512;
    10'd92: brom_out <= 64'd3324417521285869935;
    10'd348: brom_out <= 64'd4322711149969805068;
    10'd220: brom_out <= 64'd6160499120912117934;
    10'd476: brom_out <= 64'd8371723383654335520;
    10'd60: brom_out <= 64'd3866632472152804465;
    10'd316: brom_out <= 64'd5545686084666219710;
    10'd188: brom_out <= 64'd3633365094721677201;
    10'd444: brom_out <= 64'd6181880917497703341;
    10'd124: brom_out <= 64'd5775523390321313615;
    10'd380: brom_out <= 64'd6593921752856366535;
    10'd252: brom_out <= 64'd1118592617708714057;
    10'd508: brom_out <= 64'd4130478540001382116;
    10'd2: brom_out <= 64'd9150256334426485369;
    10'd258: brom_out <= 64'd2726913976235435110;
    10'd130: brom_out <= 64'd2799537887104471251;
    10'd386: brom_out <= 64'd5742128143480654282;
    10'd66: brom_out <= 64'd4848840577486999766;
    10'd322: brom_out <= 64'd5564951036314476973;
    10'd194: brom_out <= 64'd1539629244627310107;
    10'd450: brom_out <= 64'd8551637415506572346;
    10'd34: brom_out <= 64'd5569609541362591627;
    10'd290: brom_out <= 64'd3139435852145256442;
    10'd162: brom_out <= 64'd2805030511231525764;
    10'd418: brom_out <= 64'd91987351604627050;
    10'd98: brom_out <= 64'd2519301650103661960;
    10'd354: brom_out <= 64'd2610367100111832212;
    10'd226: brom_out <= 64'd3507173358449499779;
    10'd482: brom_out <= 64'd5421197279853390596;
    10'd18: brom_out <= 64'd5411415188401616703;
    10'd274: brom_out <= 64'd806771516604876704;
    10'd146: brom_out <= 64'd8252964877799973406;
    10'd402: brom_out <= 64'd4131185556170130308;
    10'd82: brom_out <= 64'd5121098992128955161;
    10'd338: brom_out <= 64'd8838718518559474163;
    10'd210: brom_out <= 64'd4217348036314092382;
    10'd466: brom_out <= 64'd8748419681862114146;
    10'd50: brom_out <= 64'd5747717726212286166;
    10'd306: brom_out <= 64'd8431525056773163324;
    10'd178: brom_out <= 64'd8135317976049821842;
    10'd434: brom_out <= 64'd3758573853795653427;
    10'd114: brom_out <= 64'd5108575401283476645;
    10'd370: brom_out <= 64'd6283534932199547339;
    10'd242: brom_out <= 64'd4633933436842356737;
    10'd498: brom_out <= 64'd911760100456784026;
    10'd10: brom_out <= 64'd6588969549873072984;
    10'd266: brom_out <= 64'd7537176118984402773;
    10'd138: brom_out <= 64'd4765782474432323605;
    10'd394: brom_out <= 64'd4784055077466289542;
    10'd74: brom_out <= 64'd695669619354178199;
    10'd330: brom_out <= 64'd3148801124557623449;
    10'd202: brom_out <= 64'd6519885780090122409;
    10'd458: brom_out <= 64'd7450817543983322844;
    10'd42: brom_out <= 64'd7396774219033937672;
    10'd298: brom_out <= 64'd5992435799082823388;
    10'd170: brom_out <= 64'd1415882188212200225;
    10'd426: brom_out <= 64'd820027634638271577;
    10'd106: brom_out <= 64'd6938251047297990533;
    10'd362: brom_out <= 64'd8673620925411977753;
    10'd234: brom_out <= 64'd1992283337758212979;
    10'd490: brom_out <= 64'd6319980041019054251;
    10'd26: brom_out <= 64'd3851039626226392450;
    10'd282: brom_out <= 64'd5711684474143641757;
    10'd154: brom_out <= 64'd6768544696756439421;
    10'd410: brom_out <= 64'd4677673593772524828;
    10'd90: brom_out <= 64'd6185725345812273456;
    10'd346: brom_out <= 64'd8312556079981528030;
    10'd218: brom_out <= 64'd8948912045682648319;
    10'd474: brom_out <= 64'd1414658525045134853;
    10'd58: brom_out <= 64'd4057166001169818856;
    10'd314: brom_out <= 64'd672919549451933827;
    10'd186: brom_out <= 64'd196307236251518595;
    10'd442: brom_out <= 64'd3445970765661623385;
    10'd122: brom_out <= 64'd6590112200699224071;
    10'd378: brom_out <= 64'd8440836487301065001;
    10'd250: brom_out <= 64'd3633265221550976288;
    10'd506: brom_out <= 64'd830325714398867404;
    10'd6: brom_out <= 64'd3293074636399430213;
    10'd262: brom_out <= 64'd9206702681534441482;
    10'd134: brom_out <= 64'd7698250944354989161;
    10'd390: brom_out <= 64'd6913663135607926584;
    10'd70: brom_out <= 64'd2862891865227566885;
    10'd326: brom_out <= 64'd5318448438505440257;
    10'd198: brom_out <= 64'd5215707159989682948;
    10'd454: brom_out <= 64'd2408543357995828304;
    10'd38: brom_out <= 64'd1331680507007219705;
    10'd294: brom_out <= 64'd789422816571225780;
    10'd166: brom_out <= 64'd1512800906605612428;
    10'd422: brom_out <= 64'd725251043603134492;
    10'd102: brom_out <= 64'd3241756220799506222;
    10'd358: brom_out <= 64'd7892653319965062638;
    10'd230: brom_out <= 64'd1144176920185415535;
    10'd486: brom_out <= 64'd6062993788722341892;
    10'd22: brom_out <= 64'd7586867602903602858;
    10'd278: brom_out <= 64'd5757481406149589238;
    10'd150: brom_out <= 64'd2703396381905810774;
    10'd406: brom_out <= 64'd5769552562384596599;
    10'd86: brom_out <= 64'd3018928514936204385;
    10'd342: brom_out <= 64'd4397702267799328608;
    10'd214: brom_out <= 64'd6481798364871042424;
    10'd470: brom_out <= 64'd3482983880212475854;
    10'd54: brom_out <= 64'd880050980480071141;
    10'd310: brom_out <= 64'd3281923340519708537;
    10'd182: brom_out <= 64'd4519341334859734073;
    10'd438: brom_out <= 64'd1337980060505609637;
    10'd118: brom_out <= 64'd8162841956676165738;
    10'd374: brom_out <= 64'd8694371873892844208;
    10'd246: brom_out <= 64'd3936667969893923919;
    10'd502: brom_out <= 64'd713405409942497823;
    10'd14: brom_out <= 64'd4290018412507268451;
    10'd270: brom_out <= 64'd1100339483998246003;
    10'd142: brom_out <= 64'd8105253848644364450;
    10'd398: brom_out <= 64'd7286314464983170863;
    10'd78: brom_out <= 64'd7530083780768442237;
    10'd334: brom_out <= 64'd4613903798598080436;
    10'd206: brom_out <= 64'd1503390632805335282;
    10'd462: brom_out <= 64'd5708860785940369427;
    10'd46: brom_out <= 64'd118243567567768095;
    10'd302: brom_out <= 64'd7077564256689660660;
    10'd174: brom_out <= 64'd1689924925158498949;
    10'd430: brom_out <= 64'd2003304190459111066;
    10'd110: brom_out <= 64'd3754010688254048597;
    10'd366: brom_out <= 64'd8513076200388136183;
    10'd238: brom_out <= 64'd3343459330700479572;
    10'd494: brom_out <= 64'd2497038050456785463;
    10'd30: brom_out <= 64'd4110036900460384796;
    10'd286: brom_out <= 64'd6501664496823873080;
    10'd158: brom_out <= 64'd6326125611953081505;
    10'd414: brom_out <= 64'd7183585907134239486;
    10'd94: brom_out <= 64'd1960716502804548672;
    10'd350: brom_out <= 64'd1985994961055839280;
    10'd222: brom_out <= 64'd3651142297411659187;
    10'd478: brom_out <= 64'd2072885801364544572;
    10'd62: brom_out <= 64'd1468430662791236228;
    10'd318: brom_out <= 64'd1435120993511282705;
    10'd190: brom_out <= 64'd5917399405983790504;
    10'd446: brom_out <= 64'd1950822828069733729;
    10'd126: brom_out <= 64'd9097630694651455464;
    10'd382: brom_out <= 64'd7427050020511569441;
    10'd254: brom_out <= 64'd8063678981840380015;
    10'd510: brom_out <= 64'd3031303078308718036;
    10'd1: brom_out <= 64'd3127052517479868225;
    10'd257: brom_out <= 64'd6914660438246835908;
    10'd129: brom_out <= 64'd8927943298820454076;
    10'd385: brom_out <= 64'd3854526127297200834;
    10'd65: brom_out <= 64'd4304180803912282259;
    10'd321: brom_out <= 64'd3119079411128405209;
    10'd193: brom_out <= 64'd7817367043308214467;
    10'd449: brom_out <= 64'd2126660867906687864;
    10'd33: brom_out <= 64'd6475240946856553091;
    10'd289: brom_out <= 64'd3032208211650146388;
    10'd161: brom_out <= 64'd9004572314107590138;
    10'd417: brom_out <= 64'd4725094368207763061;
    10'd97: brom_out <= 64'd6446311831687328438;
    10'd353: brom_out <= 64'd1478979661686592040;
    10'd225: brom_out <= 64'd8566281893646113;
    10'd481: brom_out <= 64'd333801395018402419;
    10'd17: brom_out <= 64'd1467033842096743702;
    10'd273: brom_out <= 64'd4751890286330071625;
    10'd145: brom_out <= 64'd7747822092528642924;
    10'd401: brom_out <= 64'd2777986735042830839;
    10'd81: brom_out <= 64'd8395034085139528506;
    10'd337: brom_out <= 64'd7441158198174016671;
    10'd209: brom_out <= 64'd17521832455993642;
    10'd465: brom_out <= 64'd5745260692505968145;
    10'd49: brom_out <= 64'd2943321537520600659;
    10'd305: brom_out <= 64'd6579678929095156593;
    10'd177: brom_out <= 64'd7687396513344217400;
    10'd433: brom_out <= 64'd5651215856363377316;
    10'd113: brom_out <= 64'd494499881005363032;
    10'd369: brom_out <= 64'd7462328687096900295;
    10'd241: brom_out <= 64'd1707361404853655714;
    10'd497: brom_out <= 64'd3506647722126204218;
    10'd9: brom_out <= 64'd2567313654253520317;
    10'd265: brom_out <= 64'd1778468342386166084;
    10'd137: brom_out <= 64'd2868266086180312958;
    10'd393: brom_out <= 64'd3580819943894297764;
    10'd73: brom_out <= 64'd2004505146951275140;
    10'd329: brom_out <= 64'd1737665055851572803;
    10'd201: brom_out <= 64'd4446551631123665655;
    10'd457: brom_out <= 64'd2840283348677403338;
    10'd41: brom_out <= 64'd7920402332462387511;
    10'd297: brom_out <= 64'd7125835522680848670;
    10'd169: brom_out <= 64'd3823809497424801247;
    10'd425: brom_out <= 64'd4077815017758764724;
    10'd105: brom_out <= 64'd3042490808619695370;
    10'd361: brom_out <= 64'd8341925111666110475;
    10'd233: brom_out <= 64'd1901574174662490027;
    10'd489: brom_out <= 64'd8165494333656525134;
    10'd25: brom_out <= 64'd1215003878949612048;
    10'd281: brom_out <= 64'd5269356158780504864;
    10'd153: brom_out <= 64'd8765870513679473211;
    10'd409: brom_out <= 64'd6319435406754674390;
    10'd89: brom_out <= 64'd4752592209480917425;
    10'd345: brom_out <= 64'd2931018764400806070;
    10'd217: brom_out <= 64'd962867634407305569;
    10'd473: brom_out <= 64'd8680510475920407927;
    10'd57: brom_out <= 64'd4151717614504932492;
    10'd313: brom_out <= 64'd2212864360945965123;
    10'd185: brom_out <= 64'd7149484177775971227;
    10'd441: brom_out <= 64'd8698260697543325537;
    10'd121: brom_out <= 64'd6520183508896026597;
    10'd377: brom_out <= 64'd9129774312610320619;
    10'd249: brom_out <= 64'd9123574294358671657;
    10'd505: brom_out <= 64'd2133757072145401712;
    10'd5: brom_out <= 64'd7153207102067290344;
    10'd261: brom_out <= 64'd7160540774931803866;
    10'd133: brom_out <= 64'd5541375517500192895;
    10'd389: brom_out <= 64'd4175560118002252921;
    10'd69: brom_out <= 64'd4091222591604623441;
    10'd325: brom_out <= 64'd8580562440646539131;
    10'd197: brom_out <= 64'd7055503816228831091;
    10'd453: brom_out <= 64'd4971028798941293784;
    10'd37: brom_out <= 64'd9036614214691043214;
    10'd293: brom_out <= 64'd5041872014433074100;
    10'd165: brom_out <= 64'd6265810223453665551;
    10'd421: brom_out <= 64'd3005741243809146285;
    10'd101: brom_out <= 64'd5458238346969861276;
    10'd357: brom_out <= 64'd7976876523254192230;
    10'd229: brom_out <= 64'd7990560214861353583;
    10'd485: brom_out <= 64'd2351202851047628420;
    10'd21: brom_out <= 64'd6891504871357446422;
    10'd277: brom_out <= 64'd5069629123053312106;
    10'd149: brom_out <= 64'd2857441601682776678;
    10'd405: brom_out <= 64'd8907923421314590115;
    10'd85: brom_out <= 64'd8037258735659770483;
    10'd341: brom_out <= 64'd3682273990606439039;
    10'd213: brom_out <= 64'd5880920423784685274;
    10'd469: brom_out <= 64'd9052054262515000354;
    10'd53: brom_out <= 64'd7783606212229745263;
    10'd309: brom_out <= 64'd5515184158531911546;
    10'd181: brom_out <= 64'd8240076708661524496;
    10'd437: brom_out <= 64'd5168690797098687629;
    10'd117: brom_out <= 64'd3877069780779427166;
    10'd373: brom_out <= 64'd8969075915070151768;
    10'd245: brom_out <= 64'd8632467951852587989;
    10'd501: brom_out <= 64'd7857926944957203380;
    10'd13: brom_out <= 64'd1287674294028378649;
    10'd269: brom_out <= 64'd8373705960209865750;
    10'd141: brom_out <= 64'd5410674334166473286;
    10'd397: brom_out <= 64'd4401819749409430491;
    10'd77: brom_out <= 64'd4174433604295068968;
    10'd333: brom_out <= 64'd4196968460687196785;
    10'd205: brom_out <= 64'd5852786553912777685;
    10'd461: brom_out <= 64'd4538780524597464161;
    10'd45: brom_out <= 64'd5698207036020272794;
    10'd301: brom_out <= 64'd287090937624021185;
    10'd173: brom_out <= 64'd7704688953664041795;
    10'd429: brom_out <= 64'd546478178973529773;
    10'd109: brom_out <= 64'd9168100354083393324;
    10'd365: brom_out <= 64'd6230035500739914156;
    10'd237: brom_out <= 64'd3287964157657373940;
    10'd493: brom_out <= 64'd3289458284692175700;
    10'd29: brom_out <= 64'd1821424608084578998;
    10'd285: brom_out <= 64'd6524722060171723622;
    10'd157: brom_out <= 64'd7524025148374291789;
    10'd413: brom_out <= 64'd2170069437537526133;
    10'd93: brom_out <= 64'd8528027318223251457;
    10'd349: brom_out <= 64'd6079977503648451335;
    10'd221: brom_out <= 64'd6552355050471698204;
    10'd477: brom_out <= 64'd8219861536954301229;
    10'd61: brom_out <= 64'd3063481684957609078;
    10'd317: brom_out <= 64'd1330381704714286085;
    10'd189: brom_out <= 64'd4041634879120597886;
    10'd445: brom_out <= 64'd7253780654183843384;
    10'd125: brom_out <= 64'd3651945852037892795;
    10'd381: brom_out <= 64'd3784018163499518601;
    10'd253: brom_out <= 64'd3794573246885287845;
    10'd509: brom_out <= 64'd2997007021939187347;
    10'd3: brom_out <= 64'd6825597430088558793;
    10'd259: brom_out <= 64'd4148280298264435145;
    10'd131: brom_out <= 64'd2187018093810691720;
    10'd387: brom_out <= 64'd822715829145346347;
    10'd67: brom_out <= 64'd6083010805285052716;
    10'd323: brom_out <= 64'd3036875632463858834;
    10'd195: brom_out <= 64'd2456301622261705551;
    10'd451: brom_out <= 64'd1435047781493708974;
    10'd35: brom_out <= 64'd3495906847793555496;
    10'd291: brom_out <= 64'd6846824846681755777;
    10'd163: brom_out <= 64'd4806777613109574958;
    10'd419: brom_out <= 64'd7767226473893413332;
    10'd99: brom_out <= 64'd3412151563337741352;
    10'd355: brom_out <= 64'd3368411057424669635;
    10'd227: brom_out <= 64'd6295273620685999449;
    10'd483: brom_out <= 64'd7292703967224865486;
    10'd19: brom_out <= 64'd8367416970837404480;
    10'd275: brom_out <= 64'd6060747830154195747;
    10'd147: brom_out <= 64'd1481999355516963175;
    10'd403: brom_out <= 64'd2051836413390839457;
    10'd83: brom_out <= 64'd5160625525529957528;
    10'd339: brom_out <= 64'd3854484312171404456;
    10'd211: brom_out <= 64'd2051998054788366270;
    10'd467: brom_out <= 64'd1674345919730951813;
    10'd51: brom_out <= 64'd4614122134803297477;
    10'd307: brom_out <= 64'd25054386228368260;
    10'd179: brom_out <= 64'd5991839321352371775;
    10'd435: brom_out <= 64'd6760985867545539242;
    10'd115: brom_out <= 64'd2151578802008365031;
    10'd371: brom_out <= 64'd6628447066861725489;
    10'd243: brom_out <= 64'd6447223936141958870;
    10'd499: brom_out <= 64'd4628098658155976042;
    10'd11: brom_out <= 64'd7820318430984191122;
    10'd267: brom_out <= 64'd7664280676247221904;
    10'd139: brom_out <= 64'd4633112736508198766;
    10'd395: brom_out <= 64'd4419790281338715805;
    10'd75: brom_out <= 64'd1189038338221773258;
    10'd331: brom_out <= 64'd1113248537812598346;
    10'd203: brom_out <= 64'd2086211756656440867;
    10'd459: brom_out <= 64'd6363705655307338806;
    10'd43: brom_out <= 64'd1188483528343374386;
    10'd299: brom_out <= 64'd176563187302484685;
    10'd171: brom_out <= 64'd5300966512209250050;
    10'd427: brom_out <= 64'd2595667101902401433;
    10'd107: brom_out <= 64'd6526255316566008010;
    10'd363: brom_out <= 64'd2847404267546166357;
    10'd235: brom_out <= 64'd2875223919672073068;
    10'd491: brom_out <= 64'd5252122029312962963;
    10'd27: brom_out <= 64'd6004430279489338680;
    10'd283: brom_out <= 64'd8871767897380268353;
    10'd155: brom_out <= 64'd8658919390669651664;
    10'd411: brom_out <= 64'd5511461520034253554;
    10'd91: brom_out <= 64'd4798463378767722612;
    10'd347: brom_out <= 64'd585096259269936048;
    10'd219: brom_out <= 64'd6259526245218962991;
    10'd475: brom_out <= 64'd486400348447004409;
    10'd59: brom_out <= 64'd5295131112655049137;
    10'd315: brom_out <= 64'd6072046178105556475;
    10'd187: brom_out <= 64'd1364531386125093388;
    10'd443: brom_out <= 64'd1664928300054969876;
    10'd123: brom_out <= 64'd4635191165656492150;
    10'd379: brom_out <= 64'd1755068967933061315;
    10'd251: brom_out <= 64'd6244689180377020923;
    10'd507: brom_out <= 64'd8758553949588800273;
    10'd7: brom_out <= 64'd5112583091541522973;
    10'd263: brom_out <= 64'd7835211644950567469;
    10'd135: brom_out <= 64'd5401614836719703272;
    10'd391: brom_out <= 64'd2228552985412019277;
    10'd71: brom_out <= 64'd4822434129781452362;
    10'd327: brom_out <= 64'd1078913570171309648;
    10'd199: brom_out <= 64'd5359119263554810248;
    10'd455: brom_out <= 64'd6781627562122407399;
    10'd39: brom_out <= 64'd8944063972887106670;
    10'd295: brom_out <= 64'd4822808530417619233;
    10'd167: brom_out <= 64'd4414284518212157732;
    10'd423: brom_out <= 64'd5450767261026876886;
    10'd103: brom_out <= 64'd8021309328199436730;
    10'd359: brom_out <= 64'd6199672516180526071;
    10'd231: brom_out <= 64'd2608525535082964773;
    10'd487: brom_out <= 64'd599730283692523374;
    10'd23: brom_out <= 64'd7058677087284092182;
    10'd279: brom_out <= 64'd812235029203875617;
    10'd151: brom_out <= 64'd6034460869506398985;
    10'd407: brom_out <= 64'd8947667063148711049;
    10'd87: brom_out <= 64'd1585371721068583241;
    10'd343: brom_out <= 64'd3433509905416311683;
    10'd215: brom_out <= 64'd1168596851321766456;
    10'd471: brom_out <= 64'd5032214272686406166;
    10'd55: brom_out <= 64'd5314247580215590840;
    10'd311: brom_out <= 64'd3591529433803820433;
    10'd183: brom_out <= 64'd6353718731862795407;
    10'd439: brom_out <= 64'd6411251051681906994;
    10'd119: brom_out <= 64'd1123132456013002459;
    10'd375: brom_out <= 64'd7030554445186196665;
    10'd247: brom_out <= 64'd168302224660410828;
    10'd503: brom_out <= 64'd333363560357025169;
    10'd15: brom_out <= 64'd8710174058585331351;
    10'd271: brom_out <= 64'd849306692269551679;
    10'd143: brom_out <= 64'd2464563482745670645;
    10'd399: brom_out <= 64'd9151515973652221402;
    10'd79: brom_out <= 64'd7697402264257745017;
    10'd335: brom_out <= 64'd3504473931275065124;
    10'd207: brom_out <= 64'd8759164961417563512;
    10'd463: brom_out <= 64'd6716916671807146392;
    10'd47: brom_out <= 64'd4486934250525894693;
    10'd303: brom_out <= 64'd2749009972353655762;
    10'd175: brom_out <= 64'd6919778738676338510;
    10'd431: brom_out <= 64'd3404093846247594996;
    10'd111: brom_out <= 64'd1722163249877292090;
    10'd367: brom_out <= 64'd1141842582310077908;
    10'd239: brom_out <= 64'd6889879677402930206;
    10'd495: brom_out <= 64'd7848005646647114461;
    10'd31: brom_out <= 64'd1547693224024900634;
    10'd287: brom_out <= 64'd6382089802135409144;
    10'd159: brom_out <= 64'd6658739335726264481;
    10'd415: brom_out <= 64'd4955822627172985255;
    10'd95: brom_out <= 64'd2293080637268173952;
    10'd351: brom_out <= 64'd6769971139694742693;
    10'd223: brom_out <= 64'd801305510105442737;
    10'd479: brom_out <= 64'd9096591304164137574;
    10'd63: brom_out <= 64'd1396316958451531348;
    10'd319: brom_out <= 64'd6585546512385483974;
    10'd191: brom_out <= 64'd7094683365482870580;
    10'd447: brom_out <= 64'd8631772682564570593;
    10'd127: brom_out <= 64'd8074623464407446434;
    10'd383: brom_out <= 64'd7692930341342185952;
    10'd255: brom_out <= 64'd7920910159561005345;
    10'd511: brom_out <= 64'd4803548634770013292;
    default: brom_out <= 64'h1;
    endcase
end

generate
    if(DELAY == 1) begin
        assign b = brom_out;
    end
endgenerate

endmodule

//-------------------------------------------------------------------------------------------------

module tw_rom_10_ntt_nwc
#(
    parameter LOGN  = 10,
    parameter LOGQ  = 64,
    parameter DELAY = 1,
    parameter STAGE = 10
)(
    input            clk,
    input [LOGN-1:0] raddr,
    output[LOGQ-1:0] b
);

(* ram_style = "block" *)
reg [LOGQ-1:0] brom_out, brom_out2;

always @(posedge clk) begin
    case(raddr[STAGE-1:0])
    11'd0: brom_out <= 64'd1102913100553729005;
    11'd512: brom_out <= 64'd4595731803495303327;
    11'd256: brom_out <= 64'd4005117716490349010;
    11'd768: brom_out <= 64'd2678065129254935256;
    11'd128: brom_out <= 64'd2801867022993033546;
    11'd640: brom_out <= 64'd3256237472906815544;
    11'd384: brom_out <= 64'd78521125945926901;
    11'd896: brom_out <= 64'd62383298268607752;
    11'd64: brom_out <= 64'd2038520525822259048;
    11'd576: brom_out <= 64'd8061736108804448278;
    11'd320: brom_out <= 64'd3633979900330440892;
    11'd832: brom_out <= 64'd4114200839665517402;
    11'd192: brom_out <= 64'd7574768217639654355;
    11'd704: brom_out <= 64'd8816500119098547526;
    11'd448: brom_out <= 64'd1514057220951852292;
    11'd960: brom_out <= 64'd3917320098766147730;
    11'd32: brom_out <= 64'd3702518847184112432;
    11'd544: brom_out <= 64'd8400965878765427026;
    11'd288: brom_out <= 64'd1292420980917360603;
    11'd800: brom_out <= 64'd5959304096792569751;
    11'd160: brom_out <= 64'd4369822744919577129;
    11'd672: brom_out <= 64'd8058518244289887562;
    11'd416: brom_out <= 64'd3950582044138852963;
    11'd928: brom_out <= 64'd9129940191982502832;
    11'd96: brom_out <= 64'd1189672448575511328;
    11'd608: brom_out <= 64'd6265146028599173595;
    11'd352: brom_out <= 64'd4912519834823704407;
    11'd864: brom_out <= 64'd6400216294734455669;
    11'd224: brom_out <= 64'd1203939852511973662;
    11'd736: brom_out <= 64'd6333478367606839407;
    11'd480: brom_out <= 64'd7222535658536760892;
    11'd992: brom_out <= 64'd4564125134977115371;
    11'd16: brom_out <= 64'd344548888781770986;
    11'd528: brom_out <= 64'd5218202542817394251;
    11'd272: brom_out <= 64'd335350576825950082;
    11'd784: brom_out <= 64'd3388698090164268880;
    11'd144: brom_out <= 64'd4414035617291553258;
    11'd656: brom_out <= 64'd4346661030238530214;
    11'd400: brom_out <= 64'd6162069774348355978;
    11'd912: brom_out <= 64'd905080829528335056;
    11'd80: brom_out <= 64'd5945019363494978713;
    11'd592: brom_out <= 64'd8830493778383512291;
    11'd336: brom_out <= 64'd478119158814609466;
    11'd848: brom_out <= 64'd6215685832894845107;
    11'd208: brom_out <= 64'd4215582806609882491;
    11'd720: brom_out <= 64'd3763494781935998767;
    11'd464: brom_out <= 64'd4024235301766674686;
    11'd976: brom_out <= 64'd6261499129228396190;
    11'd48: brom_out <= 64'd5160493589408218780;
    11'd560: brom_out <= 64'd6296175845735511856;
    11'd304: brom_out <= 64'd6596423659328983517;
    11'd816: brom_out <= 64'd9099378341091656482;
    11'd176: brom_out <= 64'd3827692355908478929;
    11'd688: brom_out <= 64'd3512444620723338488;
    11'd432: brom_out <= 64'd8932324166801541824;
    11'd944: brom_out <= 64'd3530957463225895281;
    11'd112: brom_out <= 64'd7500931859087234329;
    11'd624: brom_out <= 64'd6205084145235084221;
    11'd368: brom_out <= 64'd3780203902726182378;
    11'd880: brom_out <= 64'd4849251867203539042;
    11'd240: brom_out <= 64'd1121104267230146280;
    11'd752: brom_out <= 64'd1885864751055057353;
    11'd496: brom_out <= 64'd4011863120442953560;
    11'd1008: brom_out <= 64'd4797402059262399444;
    11'd8: brom_out <= 64'd7325184581455921607;
    11'd520: brom_out <= 64'd164674200546607604;
    11'd264: brom_out <= 64'd2173064029340428803;
    11'd776: brom_out <= 64'd7922160522628872772;
    11'd136: brom_out <= 64'd1779228674047657867;
    11'd648: brom_out <= 64'd8897863336940776164;
    11'd392: brom_out <= 64'd25138778867551862;
    11'd904: brom_out <= 64'd7679327987615867679;
    11'd72: brom_out <= 64'd418688512246794328;
    11'd584: brom_out <= 64'd4886014524849036326;
    11'd328: brom_out <= 64'd7670512215868297688;
    11'd840: brom_out <= 64'd3393684384123953368;
    11'd200: brom_out <= 64'd7248112848643534511;
    11'd712: brom_out <= 64'd9161163982018377625;
    11'd456: brom_out <= 64'd3183672025538269624;
    11'd968: brom_out <= 64'd7914039759715212288;
    11'd40: brom_out <= 64'd7849000344767537809;
    11'd552: brom_out <= 64'd5138973604269881666;
    11'd296: brom_out <= 64'd8374712657994971746;
    11'd808: brom_out <= 64'd6515807241519471828;
    11'd168: brom_out <= 64'd1331624447098205033;
    11'd680: brom_out <= 64'd7011739122720262005;
    11'd424: brom_out <= 64'd4802317643994205088;
    11'd936: brom_out <= 64'd5954414081382772179;
    11'd104: brom_out <= 64'd3900996048308082675;
    11'd616: brom_out <= 64'd3500901095250623076;
    11'd360: brom_out <= 64'd7605970516342646990;
    11'd872: brom_out <= 64'd8029507220670853362;
    11'd232: brom_out <= 64'd2432010159645715397;
    11'd744: brom_out <= 64'd7692433165927744565;
    11'd488: brom_out <= 64'd4082435061276421983;
    11'd1000: brom_out <= 64'd418379368903778945;
    11'd24: brom_out <= 64'd3839782310825792117;
    11'd536: brom_out <= 64'd3161833067360455250;
    11'd280: brom_out <= 64'd4777872077056980363;
    11'd792: brom_out <= 64'd5322751941608048097;
    11'd152: brom_out <= 64'd8988022062613589533;
    11'd664: brom_out <= 64'd8155382693858119578;
    11'd408: brom_out <= 64'd5693674981823269218;
    11'd920: brom_out <= 64'd7838092352335735356;
    11'd88: brom_out <= 64'd6432855811330329932;
    11'd600: brom_out <= 64'd5258779288804072394;
    11'd344: brom_out <= 64'd7660349318066984762;
    11'd856: brom_out <= 64'd5171475373150897937;
    11'd216: brom_out <= 64'd5738954251284061668;
    11'd728: brom_out <= 64'd1314283965644365680;
    11'd472: brom_out <= 64'd1083320007172303764;
    11'd984: brom_out <= 64'd8416441445159376236;
    11'd56: brom_out <= 64'd453811032764871892;
    11'd568: brom_out <= 64'd2206364998037189985;
    11'd312: brom_out <= 64'd5044057647806587586;
    11'd824: brom_out <= 64'd1745036897308546683;
    11'd184: brom_out <= 64'd1352173756344525495;
    11'd696: brom_out <= 64'd962407481846958591;
    11'd440: brom_out <= 64'd5896964627131169131;
    11'd952: brom_out <= 64'd114955450999687352;
    11'd120: brom_out <= 64'd7103911473611199541;
    11'd632: brom_out <= 64'd5549144129026746013;
    11'd376: brom_out <= 64'd9051064044881936071;
    11'd888: brom_out <= 64'd1892659099199940448;
    11'd248: brom_out <= 64'd2137770580285350027;
    11'd760: brom_out <= 64'd3707251717625885791;
    11'd504: brom_out <= 64'd6989967860725554358;
    11'd1016: brom_out <= 64'd5799824691966670023;
    11'd4: brom_out <= 64'd5667686056105230206;
    11'd516: brom_out <= 64'd1938270965119171169;
    11'd260: brom_out <= 64'd625448301026631026;
    11'd772: brom_out <= 64'd2164118330631263854;
    11'd132: brom_out <= 64'd7303964566607951423;
    11'd644: brom_out <= 64'd2310560732345386485;
    11'd388: brom_out <= 64'd402155676505531812;
    11'd900: brom_out <= 64'd7741423298594687150;
    11'd68: brom_out <= 64'd1625945569422476240;
    11'd580: brom_out <= 64'd1873889101993027220;
    11'd324: brom_out <= 64'd1313331331708123806;
    11'd836: brom_out <= 64'd5792180516837140858;
    11'd196: brom_out <= 64'd1687881817758787752;
    11'd708: brom_out <= 64'd6566502495667702930;
    11'd452: brom_out <= 64'd502463928244531822;
    11'd964: brom_out <= 64'd2080550169979121770;
    11'd36: brom_out <= 64'd819099372979029972;
    11'd548: brom_out <= 64'd2270794757509049429;
    11'd292: brom_out <= 64'd3048930568431300260;
    11'd804: brom_out <= 64'd716419806412526384;
    11'd164: brom_out <= 64'd4100239665487453604;
    11'd676: brom_out <= 64'd7417372571204481830;
    11'd420: brom_out <= 64'd7169512332837823604;
    11'd932: brom_out <= 64'd902885216720223210;
    11'd100: brom_out <= 64'd2916236583736325519;
    11'd612: brom_out <= 64'd3102877355736081607;
    11'd356: brom_out <= 64'd2158981712364655228;
    11'd868: brom_out <= 64'd8234108938174010322;
    11'd228: brom_out <= 64'd4875826095999072140;
    11'd740: brom_out <= 64'd623780653727302203;
    11'd484: brom_out <= 64'd4852120695248117336;
    11'd996: brom_out <= 64'd4782115157531486230;
    11'd20: brom_out <= 64'd3777600355184077437;
    11'd532: brom_out <= 64'd1556515623451888075;
    11'd276: brom_out <= 64'd7183671453211506471;
    11'd788: brom_out <= 64'd5028445509124063333;
    11'd148: brom_out <= 64'd3773506948494418480;
    11'd660: brom_out <= 64'd593907935894979160;
    11'd404: brom_out <= 64'd1368828974385072222;
    11'd916: brom_out <= 64'd8398591941514173618;
    11'd84: brom_out <= 64'd328762820884200268;
    11'd596: brom_out <= 64'd2193863277718000910;
    11'd340: brom_out <= 64'd7584921381365002484;
    11'd852: brom_out <= 64'd9019792797984103029;
    11'd212: brom_out <= 64'd2602683653691326026;
    11'd724: brom_out <= 64'd7445483466275733942;
    11'd468: brom_out <= 64'd8852578436638496032;
    11'd980: brom_out <= 64'd6522691292269812797;
    11'd52: brom_out <= 64'd1857577982111137819;
    11'd564: brom_out <= 64'd761655569867782735;
    11'd308: brom_out <= 64'd9102526443833176819;
    11'd820: brom_out <= 64'd9178637669322844693;
    11'd180: brom_out <= 64'd3147501462716504700;
    11'd692: brom_out <= 64'd3962315922150850049;
    11'd436: brom_out <= 64'd1933497862117067950;
    11'd948: brom_out <= 64'd4565848593636494677;
    11'd116: brom_out <= 64'd7333325376921592110;
    11'd628: brom_out <= 64'd8931667155076678830;
    11'd372: brom_out <= 64'd5375557945600039679;
    11'd884: brom_out <= 64'd5508432406675787453;
    11'd244: brom_out <= 64'd2145867268931626804;
    11'd756: brom_out <= 64'd426035889455316640;
    11'd500: brom_out <= 64'd6255317374299378826;
    11'd1012: brom_out <= 64'd1920532002935580743;
    11'd12: brom_out <= 64'd6205137676891788173;
    11'd524: brom_out <= 64'd8216051810600487589;
    11'd268: brom_out <= 64'd2000665874345772028;
    11'd780: brom_out <= 64'd6798974422792108364;
    11'd140: brom_out <= 64'd3873586375647389700;
    11'd652: brom_out <= 64'd7216151128053990306;
    11'd396: brom_out <= 64'd3941823019222225634;
    11'd908: brom_out <= 64'd5876780189316004252;
    11'd76: brom_out <= 64'd8927043086982599750;
    11'd588: brom_out <= 64'd8869096447896116182;
    11'd332: brom_out <= 64'd3415602137400722566;
    11'd844: brom_out <= 64'd585382463249167719;
    11'd204: brom_out <= 64'd5105669458685259425;
    11'd716: brom_out <= 64'd8513875384724119180;
    11'd460: brom_out <= 64'd1673469281655632698;
    11'd972: brom_out <= 64'd7870565381825619063;
    11'd44: brom_out <= 64'd5281767851388166670;
    11'd556: brom_out <= 64'd5800786890988034455;
    11'd300: brom_out <= 64'd2591362338410686344;
    11'd812: brom_out <= 64'd6693195915515107207;
    11'd172: brom_out <= 64'd5844731795589899787;
    11'd684: brom_out <= 64'd6146999979043876520;
    11'd428: brom_out <= 64'd830772712952438644;
    11'd940: brom_out <= 64'd7741012073827083232;
    11'd108: brom_out <= 64'd5025424451158582242;
    11'd620: brom_out <= 64'd5084637108789426563;
    11'd364: brom_out <= 64'd6033457957159147088;
    11'd876: brom_out <= 64'd2640079237071612813;
    11'd236: brom_out <= 64'd6209342773543205362;
    11'd748: brom_out <= 64'd7005569702398285466;
    11'd492: brom_out <= 64'd1179965516540825048;
    11'd1004: brom_out <= 64'd3884405268572847662;
    11'd28: brom_out <= 64'd3169786119895682072;
    11'd540: brom_out <= 64'd1021692220188325535;
    11'd284: brom_out <= 64'd5951489724646106101;
    11'd796: brom_out <= 64'd9036507672267599775;
    11'd156: brom_out <= 64'd8580338531199479822;
    11'd668: brom_out <= 64'd5811578762429694397;
    11'd412: brom_out <= 64'd5860301030137744471;
    11'd924: brom_out <= 64'd7068377762402013418;
    11'd92: brom_out <= 64'd2387994583949301874;
    11'd604: brom_out <= 64'd1812932789727424157;
    11'd348: brom_out <= 64'd8250164011289223786;
    11'd860: brom_out <= 64'd815693730606393862;
    11'd220: brom_out <= 64'd5868434889645250855;
    11'd732: brom_out <= 64'd132458694871421557;
    11'd476: brom_out <= 64'd3617854177990257081;
    11'd988: brom_out <= 64'd6669891205375725926;
    11'd60: brom_out <= 64'd222767951529780175;
    11'd572: brom_out <= 64'd5584850174934109096;
    11'd316: brom_out <= 64'd2781981996128691817;
    11'd828: brom_out <= 64'd3186873110017313996;
    11'd188: brom_out <= 64'd6619360377626727946;
    11'd700: brom_out <= 64'd2686589714625351870;
    11'd444: brom_out <= 64'd7607391407196645499;
    11'd956: brom_out <= 64'd1328025387181652585;
    11'd124: brom_out <= 64'd7686709619505464880;
    11'd636: brom_out <= 64'd4076427909784645200;
    11'd380: brom_out <= 64'd2327416570468869961;
    11'd892: brom_out <= 64'd166849455930454591;
    11'd252: brom_out <= 64'd5051377677337681721;
    11'd764: brom_out <= 64'd1509886436569520070;
    11'd508: brom_out <= 64'd6195679539347534888;
    11'd1020: brom_out <= 64'd5090034518991737864;
    11'd2: brom_out <= 64'd331705278823141530;
    11'd514: brom_out <= 64'd1916386186435381995;
    11'd258: brom_out <= 64'd1316412973703224049;
    11'd770: brom_out <= 64'd4586326237824140186;
    11'd130: brom_out <= 64'd9125104620207024390;
    11'd642: brom_out <= 64'd3895031829224767346;
    11'd386: brom_out <= 64'd2984424569790546779;
    11'd898: brom_out <= 64'd6822997364396815932;
    11'd66: brom_out <= 64'd4507188278956917814;
    11'd578: brom_out <= 64'd7721770747228916634;
    11'd322: brom_out <= 64'd3822681420997167602;
    11'd834: brom_out <= 64'd3887545247412752285;
    11'd194: brom_out <= 64'd3050172956909809872;
    11'd706: brom_out <= 64'd6458810129696068279;
    11'd450: brom_out <= 64'd8804964526763484820;
    11'd962: brom_out <= 64'd3748546427553799479;
    11'd34: brom_out <= 64'd494274216377378736;
    11'd546: brom_out <= 64'd5351830350077338393;
    11'd290: brom_out <= 64'd7317450101610300559;
    11'd802: brom_out <= 64'd6078180130894032113;
    11'd162: brom_out <= 64'd5773608516567397090;
    11'd674: brom_out <= 64'd2432890573058181033;
    11'd418: brom_out <= 64'd4977195593406246853;
    11'd930: brom_out <= 64'd6075271958765567578;
    11'd98: brom_out <= 64'd2103746687090801379;
    11'd610: brom_out <= 64'd4675606206018073061;
    11'd354: brom_out <= 64'd484472173182833754;
    11'd866: brom_out <= 64'd5263759361851305005;
    11'd226: brom_out <= 64'd8216179491009474193;
    11'd738: brom_out <= 64'd671685460762616247;
    11'd482: brom_out <= 64'd2460547664794426212;
    11'd994: brom_out <= 64'd7074412356985759977;
    11'd18: brom_out <= 64'd8549720275696150946;
    11'd530: brom_out <= 64'd6050565049864378024;
    11'd274: brom_out <= 64'd6610019059717728193;
    11'd786: brom_out <= 64'd8954948950927174815;
    11'd146: brom_out <= 64'd339881140317908839;
    11'd658: brom_out <= 64'd5245797325928432520;
    11'd402: brom_out <= 64'd4039886054006184193;
    11'd914: brom_out <= 64'd7549827515419954059;
    11'd82: brom_out <= 64'd5227741310768365469;
    11'd594: brom_out <= 64'd4504726022688788972;
    11'd338: brom_out <= 64'd2970910451624412054;
    11'd850: brom_out <= 64'd5082200249721761243;
    11'd210: brom_out <= 64'd8527813612084473546;
    11'd722: brom_out <= 64'd7207426732065879308;
    11'd466: brom_out <= 64'd2864923865331435467;
    11'd978: brom_out <= 64'd8213543903831367261;
    11'd50: brom_out <= 64'd7970308623799195545;
    11'd562: brom_out <= 64'd1578854839664952686;
    11'd306: brom_out <= 64'd2788184500819922894;
    11'd818: brom_out <= 64'd4997739833658486655;
    11'd178: brom_out <= 64'd8471785160522617325;
    11'd690: brom_out <= 64'd8955222256909707638;
    11'd434: brom_out <= 64'd326628130286763688;
    11'd946: brom_out <= 64'd2522950735989919033;
    11'd114: brom_out <= 64'd6887711032745255742;
    11'd626: brom_out <= 64'd3516321696517407190;
    11'd370: brom_out <= 64'd984860808516397195;
    11'd882: brom_out <= 64'd2489326655436610948;
    11'd242: brom_out <= 64'd2806490387001446027;
    11'd754: brom_out <= 64'd2477351137960909314;
    11'd498: brom_out <= 64'd6321448948253248513;
    11'd1010: brom_out <= 64'd498827655396252432;
    11'd10: brom_out <= 64'd3326814094761790440;
    11'd522: brom_out <= 64'd6779561190491316855;
    11'd266: brom_out <= 64'd666647422893437467;
    11'd778: brom_out <= 64'd5058062501522262208;
    11'd138: brom_out <= 64'd4863463436130572984;
    11'd650: brom_out <= 64'd8963917332809987708;
    11'd394: brom_out <= 64'd6925859408854431027;
    11'd906: brom_out <= 64'd8402249683953484293;
    11'd74: brom_out <= 64'd4599926363795950470;
    11'd586: brom_out <= 64'd2403098808293565319;
    11'd330: brom_out <= 64'd3414624865495540060;
    11'd842: brom_out <= 64'd5238391540599559172;
    11'd202: brom_out <= 64'd2683991028645697880;
    11'd714: brom_out <= 64'd539332076438600639;
    11'd458: brom_out <= 64'd2699311646597186707;
    11'd970: brom_out <= 64'd3366966051305126938;
    11'd42: brom_out <= 64'd4416538491726633807;
    11'd554: brom_out <= 64'd259903952847149869;
    11'd298: brom_out <= 64'd7027237905526445895;
    11'd810: brom_out <= 64'd2268799027509688551;
    11'd170: brom_out <= 64'd3517922268454075034;
    11'd682: brom_out <= 64'd8942074700439913039;
    11'd426: brom_out <= 64'd1204415582446106112;
    11'd938: brom_out <= 64'd6357006725957045398;
    11'd106: brom_out <= 64'd5226018621464696967;
    11'd618: brom_out <= 64'd1656312259292181257;
    11'd362: brom_out <= 64'd1633105308011439896;
    11'd874: brom_out <= 64'd5152612501000703728;
    11'd234: brom_out <= 64'd1772931732953384017;
    11'd746: brom_out <= 64'd5867286401481316597;
    11'd490: brom_out <= 64'd2264251713198501895;
    11'd1002: brom_out <= 64'd2296722953695232321;
    11'd26: brom_out <= 64'd5069310872664059544;
    11'd538: brom_out <= 64'd3248329190411644841;
    11'd282: brom_out <= 64'd696331007242609412;
    11'd794: brom_out <= 64'd6235368745691702325;
    11'd154: brom_out <= 64'd5215432719681743341;
    11'd666: brom_out <= 64'd6814376656091464033;
    11'd410: brom_out <= 64'd4023808547623250577;
    11'd922: brom_out <= 64'd1179528608653538977;
    11'd90: brom_out <= 64'd4975661477061904853;
    11'd602: brom_out <= 64'd3885048787610312986;
    11'd346: brom_out <= 64'd8020316467693061111;
    11'd858: brom_out <= 64'd3582037561619632849;
    11'd218: brom_out <= 64'd6623537519035813176;
    11'd730: brom_out <= 64'd2991053525981376065;
    11'd474: brom_out <= 64'd4372612876602253599;
    11'd986: brom_out <= 64'd2815234299924242613;
    11'd58: brom_out <= 64'd8426041380979419904;
    11'd570: brom_out <= 64'd6548214732868127762;
    11'd314: brom_out <= 64'd5264632850253624255;
    11'd826: brom_out <= 64'd8687882850748879926;
    11'd186: brom_out <= 64'd2475140240274188043;
    11'd698: brom_out <= 64'd4231499661440202131;
    11'd442: brom_out <= 64'd6062567962812957720;
    11'd954: brom_out <= 64'd8154865951547131798;
    11'd122: brom_out <= 64'd2203451223094322762;
    11'd634: brom_out <= 64'd3733261563727931026;
    11'd378: brom_out <= 64'd1096701672734617714;
    11'd890: brom_out <= 64'd2434856672595838747;
    11'd250: brom_out <= 64'd3442823001120628633;
    11'd762: brom_out <= 64'd855970050860984344;
    11'd506: brom_out <= 64'd3793296266665166283;
    11'd1018: brom_out <= 64'd4625028499213347781;
    11'd6: brom_out <= 64'd7172243811045393643;
    11'd518: brom_out <= 64'd5349760899881279278;
    11'd262: brom_out <= 64'd5007472984365342136;
    11'd774: brom_out <= 64'd5823730381839252049;
    11'd134: brom_out <= 64'd5923984013916025162;
    11'd646: brom_out <= 64'd634583883983266145;
    11'd390: brom_out <= 64'd2108314857132696248;
    11'd902: brom_out <= 64'd7799087759160560895;
    11'd70: brom_out <= 64'd5267269215936573461;
    11'd582: brom_out <= 64'd8744139465253655004;
    11'd326: brom_out <= 64'd189106268087547237;
    11'd838: brom_out <= 64'd5679738671843934604;
    11'd198: brom_out <= 64'd998185447878790241;
    11'd710: brom_out <= 64'd5790249722416355499;
    11'd454: brom_out <= 64'd4101511390806188959;
    11'd966: brom_out <= 64'd6578345984344235708;
    11'd38: brom_out <= 64'd5208933208073689448;
    11'd550: brom_out <= 64'd8461937665451657542;
    11'd294: brom_out <= 64'd8708749152152484117;
    11'd806: brom_out <= 64'd3873551248534087511;
    11'd166: brom_out <= 64'd7157945453815143715;
    11'd678: brom_out <= 64'd8177505488046858016;
    11'd422: brom_out <= 64'd3671551594854379962;
    11'd934: brom_out <= 64'd7477596686818285089;
    11'd102: brom_out <= 64'd3520800072367565818;
    11'd614: brom_out <= 64'd4318098524395396650;
    11'd358: brom_out <= 64'd760364662072605816;
    11'd870: brom_out <= 64'd6466654536513188581;
    11'd230: brom_out <= 64'd1006312549628104935;
    11'd742: brom_out <= 64'd268999905903068517;
    11'd486: brom_out <= 64'd2544517863417907900;
    11'd998: brom_out <= 64'd6602550468570056359;
    11'd22: brom_out <= 64'd331112463124969936;
    11'd534: brom_out <= 64'd5548372674297715787;
    11'd278: brom_out <= 64'd3002431078669018093;
    11'd790: brom_out <= 64'd8614484543584024473;
    11'd150: brom_out <= 64'd7801453391915490838;
    11'd662: brom_out <= 64'd1400719953817300295;
    11'd406: brom_out <= 64'd2548864131226053734;
    11'd918: brom_out <= 64'd7186447650655557536;
    11'd86: brom_out <= 64'd2887841837436318313;
    11'd598: brom_out <= 64'd5950625068259854648;
    11'd342: brom_out <= 64'd5006322225260249573;
    11'd854: brom_out <= 64'd3901615430265803360;
    11'd214: brom_out <= 64'd8008558357275281990;
    11'd726: brom_out <= 64'd6403028868537790655;
    11'd470: brom_out <= 64'd1193634655463454607;
    11'd982: brom_out <= 64'd7901443076583028786;
    11'd54: brom_out <= 64'd7685174008941584275;
    11'd566: brom_out <= 64'd7462540017383874819;
    11'd310: brom_out <= 64'd4010273547781768614;
    11'd822: brom_out <= 64'd3024775562432476191;
    11'd182: brom_out <= 64'd8308285389689614985;
    11'd694: brom_out <= 64'd8052177048263815731;
    11'd438: brom_out <= 64'd8292868431172674679;
    11'd950: brom_out <= 64'd6710867888635545364;
    11'd118: brom_out <= 64'd765045619723753688;
    11'd630: brom_out <= 64'd5342489680170388343;
    11'd374: brom_out <= 64'd4774005550677405386;
    11'd886: brom_out <= 64'd1524367001083692685;
    11'd246: brom_out <= 64'd5209222732708414539;
    11'd758: brom_out <= 64'd2013262658437665285;
    11'd502: brom_out <= 64'd592321105965206016;
    11'd1014: brom_out <= 64'd2077143712079454508;
    11'd14: brom_out <= 64'd6624943704144324919;
    11'd526: brom_out <= 64'd8823402378843521219;
    11'd270: brom_out <= 64'd8577479475597382168;
    11'd782: brom_out <= 64'd7122058084065222170;
    11'd142: brom_out <= 64'd4899537041491779759;
    11'd654: brom_out <= 64'd8903487350221356454;
    11'd398: brom_out <= 64'd2104513439566953500;
    11'd910: brom_out <= 64'd292996083201336963;
    11'd78: brom_out <= 64'd6037508690161556393;
    11'd590: brom_out <= 64'd6531604368224188806;
    11'd334: brom_out <= 64'd7025983680737965395;
    11'd846: brom_out <= 64'd62214353023950165;
    11'd206: brom_out <= 64'd7293739831641998651;
    11'd718: brom_out <= 64'd9079580109520213237;
    11'd462: brom_out <= 64'd2714382757628886923;
    11'd974: brom_out <= 64'd4681885771850953136;
    11'd46: brom_out <= 64'd5290510743141442020;
    11'd558: brom_out <= 64'd6105427606278424468;
    11'd302: brom_out <= 64'd6735328272190945037;
    11'd814: brom_out <= 64'd3816207022314241251;
    11'd174: brom_out <= 64'd2073611639215184113;
    11'd686: brom_out <= 64'd1425902537865729979;
    11'd430: brom_out <= 64'd6640817230316013339;
    11'd942: brom_out <= 64'd2843344465769147130;
    11'd110: brom_out <= 64'd224320552559350026;
    11'd622: brom_out <= 64'd5700300283373190385;
    11'd366: brom_out <= 64'd1384350578725038654;
    11'd878: brom_out <= 64'd3482685859946588622;
    11'd238: brom_out <= 64'd2802120147652768839;
    11'd750: brom_out <= 64'd6767449512620135517;
    11'd494: brom_out <= 64'd996377262630989551;
    11'd1006: brom_out <= 64'd7094757395937096739;
    11'd30: brom_out <= 64'd7758685808708086097;
    11'd542: brom_out <= 64'd162862229894596551;
    11'd286: brom_out <= 64'd476664286229091365;
    11'd798: brom_out <= 64'd6729280471890946438;
    11'd158: brom_out <= 64'd3010982391224114088;
    11'd670: brom_out <= 64'd2958152679937921299;
    11'd414: brom_out <= 64'd5598236424952292337;
    11'd926: brom_out <= 64'd9000423794924863478;
    11'd94: brom_out <= 64'd9058002763678952859;
    11'd606: brom_out <= 64'd2520032607121689713;
    11'd350: brom_out <= 64'd7935001385118833413;
    11'd862: brom_out <= 64'd8593145202619771701;
    11'd222: brom_out <= 64'd2426069432682723438;
    11'd734: brom_out <= 64'd8501478292815056322;
    11'd478: brom_out <= 64'd23757372729667867;
    11'd990: brom_out <= 64'd6023400386987486231;
    11'd62: brom_out <= 64'd4481386419402181357;
    11'd574: brom_out <= 64'd7110429745811052508;
    11'd318: brom_out <= 64'd3023184176706965674;
    11'd830: brom_out <= 64'd8700108686837974136;
    11'd190: brom_out <= 64'd4682354897801007425;
    11'd702: brom_out <= 64'd6524547434638763383;
    11'd446: brom_out <= 64'd4337748426843001873;
    11'd958: brom_out <= 64'd2231951319336376728;
    11'd126: brom_out <= 64'd4390718853010686896;
    11'd638: brom_out <= 64'd4287893524448971608;
    11'd382: brom_out <= 64'd6751843302554367241;
    11'd894: brom_out <= 64'd7783916570026358453;
    11'd254: brom_out <= 64'd5546600636589182767;
    11'd766: brom_out <= 64'd6810071412848208525;
    11'd510: brom_out <= 64'd792070567551351799;
    11'd1022: brom_out <= 64'd3528552613765459030;
    11'd1: brom_out <= 64'd1527009950824020455;
    11'd513: brom_out <= 64'd3173670304377726411;
    11'd257: brom_out <= 64'd5166836646587597065;
    11'd769: brom_out <= 64'd1676519968667390242;
    11'd129: brom_out <= 64'd2918757492399093761;
    11'd641: brom_out <= 64'd4184126388409380134;
    11'd385: brom_out <= 64'd5823169037746669754;
    11'd897: brom_out <= 64'd7816775377648000771;
    11'd65: brom_out <= 64'd5587791659679814202;
    11'd577: brom_out <= 64'd2822778535989408567;
    11'd321: brom_out <= 64'd5832136871207562377;
    11'd833: brom_out <= 64'd3433750853083519277;
    11'd193: brom_out <= 64'd4643101887081870411;
    11'd705: brom_out <= 64'd563696475519026428;
    11'd449: brom_out <= 64'd9117853174285888050;
    11'd961: brom_out <= 64'd7220428068555961202;
    11'd33: brom_out <= 64'd5445518581501875667;
    11'd545: brom_out <= 64'd4082192015958411523;
    11'd289: brom_out <= 64'd7425855313841445797;
    11'd801: brom_out <= 64'd1809521424258670838;
    11'd161: brom_out <= 64'd7392630178923620229;
    11'd673: brom_out <= 64'd5165561524482769986;
    11'd417: brom_out <= 64'd5402496919907892894;
    11'd929: brom_out <= 64'd4390475210111465648;
    11'd97: brom_out <= 64'd4047332604529772758;
    11'd609: brom_out <= 64'd6250779680011007694;
    11'd353: brom_out <= 64'd7129037378186886574;
    11'd865: brom_out <= 64'd1319517056341783842;
    11'd225: brom_out <= 64'd6605244667463568635;
    11'd737: brom_out <= 64'd7178172838362117853;
    11'd481: brom_out <= 64'd8372383270641797411;
    11'd993: brom_out <= 64'd6822183555527485407;
    11'd17: brom_out <= 64'd1572845108645829558;
    11'd529: brom_out <= 64'd2520132840412007274;
    11'd273: brom_out <= 64'd7106724961015418341;
    11'd785: brom_out <= 64'd1292270614421363347;
    11'd145: brom_out <= 64'd1642318664855664016;
    11'd657: brom_out <= 64'd1393076932459315047;
    11'd401: brom_out <= 64'd1088076550595330003;
    11'd913: brom_out <= 64'd8024688023385731279;
    11'd81: brom_out <= 64'd4374432210238539416;
    11'd593: brom_out <= 64'd2223491687363304360;
    11'd337: brom_out <= 64'd9222684029687266857;
    11'd849: brom_out <= 64'd3709366288716809584;
    11'd209: brom_out <= 64'd8013752277862596731;
    11'd721: brom_out <= 64'd5253324035467520156;
    11'd465: brom_out <= 64'd4867650036211325578;
    11'd977: brom_out <= 64'd5357778098061340193;
    11'd49: brom_out <= 64'd2125871470203471318;
    11'd561: brom_out <= 64'd4953097448697532735;
    11'd305: brom_out <= 64'd4526467801563614800;
    11'd817: brom_out <= 64'd704204137755443298;
    11'd177: brom_out <= 64'd8381509481982198757;
    11'd689: brom_out <= 64'd6738164926973299742;
    11'd433: brom_out <= 64'd813325539083547321;
    11'd945: brom_out <= 64'd1941565973332653447;
    11'd113: brom_out <= 64'd3907478483338414094;
    11'd625: brom_out <= 64'd8880750789267131080;
    11'd369: brom_out <= 64'd6813168121181337925;
    11'd881: brom_out <= 64'd2366126602436718469;
    11'd241: brom_out <= 64'd9204011995672087541;
    11'd753: brom_out <= 64'd9081318113255327118;
    11'd497: brom_out <= 64'd5294995080171998451;
    11'd1009: brom_out <= 64'd4563606578771979378;
    11'd9: brom_out <= 64'd6682290189906599342;
    11'd521: brom_out <= 64'd6615260160847664585;
    11'd265: brom_out <= 64'd2499747760317348668;
    11'd777: brom_out <= 64'd220774408946330784;
    11'd137: brom_out <= 64'd6435347175821900655;
    11'd649: brom_out <= 64'd6643848106357390455;
    11'd393: brom_out <= 64'd6191071447783597483;
    11'd905: brom_out <= 64'd8516742478246974777;
    11'd73: brom_out <= 64'd8897437151834909042;
    11'd585: brom_out <= 64'd9032699219067860781;
    11'd329: brom_out <= 64'd1700990274694725704;
    11'd841: brom_out <= 64'd4572460370399290474;
    11'd201: brom_out <= 64'd6806940559200776408;
    11'd713: brom_out <= 64'd5562682736650988466;
    11'd457: brom_out <= 64'd4648179036277464614;
    11'd969: brom_out <= 64'd5663777043287975940;
    11'd41: brom_out <= 64'd3614648718488622517;
    11'd553: brom_out <= 64'd8025602516218589744;
    11'd297: brom_out <= 64'd5510182198338588319;
    11'd809: brom_out <= 64'd7251072921457186698;
    11'd169: brom_out <= 64'd3460988223109260373;
    11'd681: brom_out <= 64'd2855397955646245100;
    11'd425: brom_out <= 64'd8876448235781091709;
    11'd937: brom_out <= 64'd874093145357780858;
    11'd105: brom_out <= 64'd7126809288095688532;
    11'd617: brom_out <= 64'd601771167641863668;
    11'd361: brom_out <= 64'd864420952012544153;
    11'd873: brom_out <= 64'd2521421605044512323;
    11'd233: brom_out <= 64'd7521624398464494394;
    11'd745: brom_out <= 64'd8199554349178138502;
    11'd489: brom_out <= 64'd3440900081023092332;
    11'd1001: brom_out <= 64'd5116562701081850885;
    11'd25: brom_out <= 64'd6615922998039242763;
    11'd537: brom_out <= 64'd2122828736867373768;
    11'd281: brom_out <= 64'd6495472315871052654;
    11'd793: brom_out <= 64'd615834550689196678;
    11'd153: brom_out <= 64'd3496349151480100481;
    11'd665: brom_out <= 64'd4889370594359438957;
    11'd409: brom_out <= 64'd5447452542047891116;
    11'd921: brom_out <= 64'd2506350271925135261;
    11'd89: brom_out <= 64'd4625169900183292974;
    11'd601: brom_out <= 64'd3642262225836421716;
    11'd345: brom_out <= 64'd3544520116357534828;
    11'd857: brom_out <= 64'd8414575406705992960;
    11'd217: brom_out <= 64'd4059622768511913746;
    11'd729: brom_out <= 64'd468569663261293589;
    11'd473: brom_out <= 64'd456706321385894513;
    11'd985: brom_out <= 64'd8480219384681450441;
    11'd57: brom_out <= 64'd4326695183155906556;
    11'd569: brom_out <= 64'd4812882446374196222;
    11'd313: brom_out <= 64'd8355797756938721784;
    11'd825: brom_out <= 64'd7080205292498256390;
    11'd185: brom_out <= 64'd3261813778574482554;
    11'd697: brom_out <= 64'd8140874147456852453;
    11'd441: brom_out <= 64'd2167999302398932480;
    11'd953: brom_out <= 64'd7618198269109257018;
    11'd121: brom_out <= 64'd2104670626740145188;
    11'd633: brom_out <= 64'd1343223045376093288;
    11'd377: brom_out <= 64'd6303308488427599573;
    11'd889: brom_out <= 64'd1927462247068273250;
    11'd249: brom_out <= 64'd7086563346910060429;
    11'd761: brom_out <= 64'd7071548278656136848;
    11'd505: brom_out <= 64'd5653837848356806718;
    11'd1017: brom_out <= 64'd113075564764729104;
    11'd5: brom_out <= 64'd7706649108346001651;
    11'd517: brom_out <= 64'd7543858027698518528;
    11'd261: brom_out <= 64'd6139871726171298472;
    11'd773: brom_out <= 64'd4007459461997400903;
    11'd133: brom_out <= 64'd4368601964820485477;
    11'd645: brom_out <= 64'd7216537363218896285;
    11'd389: brom_out <= 64'd331508909586663393;
    11'd901: brom_out <= 64'd501434621617250977;
    11'd69: brom_out <= 64'd5345829616181158893;
    11'd581: brom_out <= 64'd3457656149741362258;
    11'd325: brom_out <= 64'd585413331536420342;
    11'd837: brom_out <= 64'd7166490740407512639;
    11'd197: brom_out <= 64'd61829322818278264;
    11'd709: brom_out <= 64'd8878323482694811936;
    11'd453: brom_out <= 64'd6797135268318975993;
    11'd965: brom_out <= 64'd3298163028476833569;
    11'd37: brom_out <= 64'd1757503418561083295;
    11'd549: brom_out <= 64'd220166632239457975;
    11'd293: brom_out <= 64'd3642980676160988416;
    11'd805: brom_out <= 64'd5182512363142578659;
    11'd165: brom_out <= 64'd6197181412830849464;
    11'd677: brom_out <= 64'd5201503226485455237;
    11'd421: brom_out <= 64'd5075818161597640077;
    11'd933: brom_out <= 64'd2940843062971874248;
    11'd101: brom_out <= 64'd7181474872531538448;
    11'd613: brom_out <= 64'd5362137396733491930;
    11'd357: brom_out <= 64'd2753317697438201979;
    11'd869: brom_out <= 64'd122506550756017413;
    11'd229: brom_out <= 64'd143958327396720651;
    11'd741: brom_out <= 64'd8163830362846381072;
    11'd485: brom_out <= 64'd587698803814343080;
    11'd997: brom_out <= 64'd4676447342981270542;
    11'd21: brom_out <= 64'd5984646794750834878;
    11'd533: brom_out <= 64'd3261485979621056498;
    11'd277: brom_out <= 64'd6926826029504761109;
    11'd789: brom_out <= 64'd6012239089180365601;
    11'd149: brom_out <= 64'd7508137942481891379;
    11'd661: brom_out <= 64'd4335064197964659539;
    11'd405: brom_out <= 64'd3515341576481069642;
    11'd917: brom_out <= 64'd1851285243088295653;
    11'd85: brom_out <= 64'd3958484914374424336;
    11'd597: brom_out <= 64'd6954783923074474543;
    11'd341: brom_out <= 64'd5070366903226930676;
    11'd853: brom_out <= 64'd2558689606074079344;
    11'd213: brom_out <= 64'd6146878404415362577;
    11'd725: brom_out <= 64'd4594800911237165801;
    11'd469: brom_out <= 64'd2784125964689156344;
    11'd981: brom_out <= 64'd8879506357919806857;
    11'd53: brom_out <= 64'd6186730927293561609;
    11'd565: brom_out <= 64'd9064173460967769874;
    11'd309: brom_out <= 64'd5187244564822774566;
    11'd821: brom_out <= 64'd5227644328066207813;
    11'd181: brom_out <= 64'd3785970388161490303;
    11'd693: brom_out <= 64'd2509718512183293069;
    11'd437: brom_out <= 64'd5758110218168465728;
    11'd949: brom_out <= 64'd4814867419846616074;
    11'd117: brom_out <= 64'd2683430372073479744;
    11'd629: brom_out <= 64'd7789650034503307067;
    11'd373: brom_out <= 64'd6807433264447476885;
    11'd885: brom_out <= 64'd4183341191108191639;
    11'd245: brom_out <= 64'd7207749336182051669;
    11'd757: brom_out <= 64'd1389138119124998720;
    11'd501: brom_out <= 64'd7385984052681800207;
    11'd1013: brom_out <= 64'd6122157121651334895;
    11'd13: brom_out <= 64'd1238696719636161094;
    11'd525: brom_out <= 64'd5981994135735259692;
    11'd269: brom_out <= 64'd516117442035369156;
    11'd781: brom_out <= 64'd4700118327586250533;
    11'd141: brom_out <= 64'd8216846839876223100;
    11'd653: brom_out <= 64'd1341898580837423017;
    11'd397: brom_out <= 64'd1649380730009983717;
    11'd909: brom_out <= 64'd4703808339260184091;
    11'd77: brom_out <= 64'd8668330478160946558;
    11'd589: brom_out <= 64'd3663232130631177082;
    11'd333: brom_out <= 64'd581076090402175181;
    11'd845: brom_out <= 64'd2221481776280657367;
    11'd205: brom_out <= 64'd5888155221788109374;
    11'd717: brom_out <= 64'd1584884239282854430;
    11'd461: brom_out <= 64'd3249217722349422785;
    11'd973: brom_out <= 64'd2017703862402965552;
    11'd45: brom_out <= 64'd4765428132147807493;
    11'd557: brom_out <= 64'd3414716947497933073;
    11'd301: brom_out <= 64'd9008273559910712642;
    11'd813: brom_out <= 64'd6757311289111676977;
    11'd173: brom_out <= 64'd4925083064398185451;
    11'd685: brom_out <= 64'd9000490380987386148;
    11'd429: brom_out <= 64'd2634628254352179088;
    11'd941: brom_out <= 64'd4946289342964105799;
    11'd109: brom_out <= 64'd3219436865258312315;
    11'd621: brom_out <= 64'd4722336290825604735;
    11'd365: brom_out <= 64'd1100322559612223103;
    11'd877: brom_out <= 64'd4740339309841169896;
    11'd237: brom_out <= 64'd2739817607316069076;
    11'd749: brom_out <= 64'd8317491426765841036;
    11'd493: brom_out <= 64'd1704950911325584250;
    11'd1005: brom_out <= 64'd3186532348549307234;
    11'd29: brom_out <= 64'd957479872005410401;
    11'd541: brom_out <= 64'd371088353612679558;
    11'd285: brom_out <= 64'd9087061851861541574;
    11'd797: brom_out <= 64'd6118620384573872227;
    11'd157: brom_out <= 64'd8594835602539730064;
    11'd669: brom_out <= 64'd1091320823777447142;
    11'd413: brom_out <= 64'd7516231720080428053;
    11'd925: brom_out <= 64'd3322253652462601701;
    11'd93: brom_out <= 64'd3670854517306604647;
    11'd605: brom_out <= 64'd8721513482441044300;
    11'd349: brom_out <= 64'd1418499548803264809;
    11'd861: brom_out <= 64'd7527660023201710545;
    11'd221: brom_out <= 64'd1345532271632170682;
    11'd733: brom_out <= 64'd917141149160099628;
    11'd477: brom_out <= 64'd2333919523156828507;
    11'd989: brom_out <= 64'd8918266820007170405;
    11'd61: brom_out <= 64'd8106152487619506999;
    11'd573: brom_out <= 64'd3805392669830113515;
    11'd317: brom_out <= 64'd5126919642324647453;
    11'd829: brom_out <= 64'd1714483633892986712;
    11'd189: brom_out <= 64'd1296572473256973960;
    11'd701: brom_out <= 64'd1882086957153388148;
    11'd445: brom_out <= 64'd6030263012495362676;
    11'd957: brom_out <= 64'd7266317117570346595;
    11'd125: brom_out <= 64'd8995510598615158165;
    11'd637: brom_out <= 64'd995086951603849713;
    11'd381: brom_out <= 64'd8636091743291140867;
    11'd893: brom_out <= 64'd1781769378676842139;
    11'd253: brom_out <= 64'd2191685270051714447;
    11'd765: brom_out <= 64'd2656374355877288154;
    11'd509: brom_out <= 64'd4987501261148305465;
    11'd1021: brom_out <= 64'd3542987084829734975;
    11'd3: brom_out <= 64'd4972921688478999892;
    11'd515: brom_out <= 64'd4784390490314142871;
    11'd259: brom_out <= 64'd6859486595377746448;
    11'd771: brom_out <= 64'd6026366267866628186;
    11'd131: brom_out <= 64'd7003030798630255435;
    11'd643: brom_out <= 64'd9155661255527747178;
    11'd387: brom_out <= 64'd2826193018771081104;
    11'd899: brom_out <= 64'd7067652521121856833;
    11'd67: brom_out <= 64'd2922269551779043038;
    11'd579: brom_out <= 64'd2295262262072788052;
    11'd323: brom_out <= 64'd13846368282169064;
    11'd835: brom_out <= 64'd270433545850009328;
    11'd195: brom_out <= 64'd39054179753570328;
    11'd707: brom_out <= 64'd3489052947642352681;
    11'd451: brom_out <= 64'd3123787049644773702;
    11'd963: brom_out <= 64'd2078333833292311636;
    11'd35: brom_out <= 64'd1476514077331314976;
    11'd547: brom_out <= 64'd542606181224160151;
    11'd291: brom_out <= 64'd8115948946013618884;
    11'd803: brom_out <= 64'd2522336249437108104;
    11'd163: brom_out <= 64'd6184511926724241706;
    11'd675: brom_out <= 64'd4040582382191874932;
    11'd419: brom_out <= 64'd1485900908579781315;
    11'd931: brom_out <= 64'd797287633007989097;
    11'd99: brom_out <= 64'd13677257000361224;
    11'd611: brom_out <= 64'd2052037289703534027;
    11'd355: brom_out <= 64'd6909328800562532699;
    11'd867: brom_out <= 64'd1839077451479082854;
    11'd227: brom_out <= 64'd3238882406020454937;
    11'd739: brom_out <= 64'd3897349523513245448;
    11'd483: brom_out <= 64'd8279003718731922783;
    11'd995: brom_out <= 64'd1094028519425961855;
    11'd19: brom_out <= 64'd9089944754788158967;
    11'd531: brom_out <= 64'd8104824511528610961;
    11'd275: brom_out <= 64'd7318335930499649148;
    11'd787: brom_out <= 64'd3288117840036850138;
    11'd147: brom_out <= 64'd6254333483692308558;
    11'd659: brom_out <= 64'd2418821237100432937;
    11'd403: brom_out <= 64'd4530139836433554292;
    11'd915: brom_out <= 64'd7970310816677404075;
    11'd83: brom_out <= 64'd2473325997743944052;
    11'd595: brom_out <= 64'd9027321022514621789;
    11'd339: brom_out <= 64'd8629179470676055812;
    11'd851: brom_out <= 64'd2646830679214791143;
    11'd211: brom_out <= 64'd7318487377759942214;
    11'd723: brom_out <= 64'd1472757774526024785;
    11'd467: brom_out <= 64'd9208255149800298927;
    11'd979: brom_out <= 64'd7997705093244106770;
    11'd51: brom_out <= 64'd6376806131588433218;
    11'd563: brom_out <= 64'd198276819140143772;
    11'd307: brom_out <= 64'd4057006210167085562;
    11'd819: brom_out <= 64'd8315450962467588491;
    11'd179: brom_out <= 64'd8890166281502929697;
    11'd691: brom_out <= 64'd6888711580551652825;
    11'd435: brom_out <= 64'd1290930582866351128;
    11'd947: brom_out <= 64'd4928029787718124417;
    11'd115: brom_out <= 64'd6460853876874714811;
    11'd627: brom_out <= 64'd3975183427385598615;
    11'd371: brom_out <= 64'd6230788417987498078;
    11'd883: brom_out <= 64'd846810251056707812;
    11'd243: brom_out <= 64'd6903342917993908620;
    11'd755: brom_out <= 64'd6552917894363667778;
    11'd499: brom_out <= 64'd3039518500019049569;
    11'd1011: brom_out <= 64'd6339147614357192038;
    11'd11: brom_out <= 64'd5020486994570292715;
    11'd523: brom_out <= 64'd6015795952029749156;
    11'd267: brom_out <= 64'd216156902476935823;
    11'd779: brom_out <= 64'd3173784488041209200;
    11'd139: brom_out <= 64'd6904042720651947488;
    11'd651: brom_out <= 64'd3047197073143512046;
    11'd395: brom_out <= 64'd2851277803142913097;
    11'd907: brom_out <= 64'd1565712890855058017;
    11'd75: brom_out <= 64'd6430137174595182183;
    11'd587: brom_out <= 64'd8647626436894153339;
    11'd331: brom_out <= 64'd4580895004721707237;
    11'd843: brom_out <= 64'd5586233649254080813;
    11'd203: brom_out <= 64'd1552474800957627860;
    11'd715: brom_out <= 64'd6277239556914161008;
    11'd459: brom_out <= 64'd8130859604558591146;
    11'd971: brom_out <= 64'd8380172696664431219;
    11'd43: brom_out <= 64'd4987120826118502355;
    11'd555: brom_out <= 64'd4014783758903962557;
    11'd299: brom_out <= 64'd3787408563903770001;
    11'd811: brom_out <= 64'd6380806961761902536;
    11'd171: brom_out <= 64'd7433176994362088473;
    11'd683: brom_out <= 64'd7528195295407567929;
    11'd427: brom_out <= 64'd6904517509735436689;
    11'd939: brom_out <= 64'd3119795926878188610;
    11'd107: brom_out <= 64'd3590495931749359103;
    11'd619: brom_out <= 64'd8012349467558720615;
    11'd363: brom_out <= 64'd1739832632716235247;
    11'd875: brom_out <= 64'd1586036392611317199;
    11'd235: brom_out <= 64'd5821703083043290091;
    11'd747: brom_out <= 64'd3137606336581079208;
    11'd491: brom_out <= 64'd3154382174460298506;
    11'd1003: brom_out <= 64'd7262846507307089798;
    11'd27: brom_out <= 64'd543826894803705978;
    11'd539: brom_out <= 64'd5096141494837811524;
    11'd283: brom_out <= 64'd6853549056042485036;
    11'd795: brom_out <= 64'd5204306756936923712;
    11'd155: brom_out <= 64'd4108995439916808286;
    11'd667: brom_out <= 64'd7707838255361434376;
    11'd411: brom_out <= 64'd6096433046458680369;
    11'd923: brom_out <= 64'd5098416780702440734;
    11'd91: brom_out <= 64'd2851129277900631036;
    11'd603: brom_out <= 64'd7277929510343960039;
    11'd347: brom_out <= 64'd2993034213610705855;
    11'd859: brom_out <= 64'd5586732638848740465;
    11'd219: brom_out <= 64'd1585427658453945272;
    11'd731: brom_out <= 64'd4841250990366375746;
    11'd475: brom_out <= 64'd3815719428901871649;
    11'd987: brom_out <= 64'd3737566005788852338;
    11'd59: brom_out <= 64'd4350436591725259429;
    11'd571: brom_out <= 64'd6200279617731237344;
    11'd315: brom_out <= 64'd1586452688103683977;
    11'd827: brom_out <= 64'd597184167161759606;
    11'd187: brom_out <= 64'd8728287108636576294;
    11'd699: brom_out <= 64'd2450795518335383150;
    11'd443: brom_out <= 64'd3864165031077615023;
    11'd955: brom_out <= 64'd6704025482711792486;
    11'd123: brom_out <= 64'd7972835908627627311;
    11'd635: brom_out <= 64'd36022640168924989;
    11'd379: brom_out <= 64'd4228600194548570995;
    11'd891: brom_out <= 64'd4643807501097303714;
    11'd251: brom_out <= 64'd968497301989212927;
    11'd763: brom_out <= 64'd8516443880759784307;
    11'd507: brom_out <= 64'd6231911985272121732;
    11'd1019: brom_out <= 64'd8461727611525100825;
    11'd7: brom_out <= 64'd3948706956136277229;
    11'd519: brom_out <= 64'd5390736926471664788;
    11'd263: brom_out <= 64'd6007025510947175156;
    11'd775: brom_out <= 64'd642913437998720848;
    11'd135: brom_out <= 64'd1194702245926272972;
    11'd647: brom_out <= 64'd2242810203672903028;
    11'd391: brom_out <= 64'd4314974606150836240;
    11'd903: brom_out <= 64'd1082513074530133782;
    11'd71: brom_out <= 64'd8152988480412639353;
    11'd583: brom_out <= 64'd1606167506240542843;
    11'd327: brom_out <= 64'd1637309547778421810;
    11'd839: brom_out <= 64'd4307950442227902464;
    11'd199: brom_out <= 64'd1014540976961417578;
    11'd711: brom_out <= 64'd3703586401268449278;
    11'd455: brom_out <= 64'd8303740360864384825;
    11'd967: brom_out <= 64'd2984492509020460139;
    11'd39: brom_out <= 64'd5002790962071147126;
    11'd551: brom_out <= 64'd6700911579012967260;
    11'd295: brom_out <= 64'd1000681170679138810;
    11'd807: brom_out <= 64'd2321442173369150588;
    11'd167: brom_out <= 64'd1656556474370501420;
    11'd679: brom_out <= 64'd2919958029833209633;
    11'd423: brom_out <= 64'd2896324170644098685;
    11'd935: brom_out <= 64'd1900135137736299752;
    11'd103: brom_out <= 64'd4254624995020049834;
    11'd615: brom_out <= 64'd608396834745710365;
    11'd359: brom_out <= 64'd3039730646554404637;
    11'd871: brom_out <= 64'd8403500667367406851;
    11'd231: brom_out <= 64'd3818591566592158579;
    11'd743: brom_out <= 64'd2439176352400363216;
    11'd487: brom_out <= 64'd6219209598344493322;
    11'd999: brom_out <= 64'd5174059410693853581;
    11'd23: brom_out <= 64'd8404649338598950687;
    11'd535: brom_out <= 64'd8163551390154089839;
    11'd279: brom_out <= 64'd5331734343637620507;
    11'd791: brom_out <= 64'd4583713786487905006;
    11'd151: brom_out <= 64'd2642030319808362412;
    11'd663: brom_out <= 64'd6536107692361147554;
    11'd407: brom_out <= 64'd1191926010696125333;
    11'd919: brom_out <= 64'd2746303970045943107;
    11'd87: brom_out <= 64'd8745925251385352737;
    11'd599: brom_out <= 64'd6714068005318992750;
    11'd343: brom_out <= 64'd1792685860936897610;
    11'd855: brom_out <= 64'd3645042965713073379;
    11'd215: brom_out <= 64'd3949377814362547728;
    11'd727: brom_out <= 64'd1519567052495348237;
    11'd471: brom_out <= 64'd4858729015412237653;
    11'd983: brom_out <= 64'd1715018151296686515;
    11'd55: brom_out <= 64'd5215512869855517538;
    11'd567: brom_out <= 64'd7580464959537686266;
    11'd311: brom_out <= 64'd8119863567815308140;
    11'd823: brom_out <= 64'd7613867444966436683;
    11'd183: brom_out <= 64'd3145699679273069605;
    11'd695: brom_out <= 64'd6044746018222371047;
    11'd439: brom_out <= 64'd1415788218295337537;
    11'd951: brom_out <= 64'd3831753525239012364;
    11'd119: brom_out <= 64'd7386813248718022410;
    11'd631: brom_out <= 64'd2905515105513391987;
    11'd375: brom_out <= 64'd4612786026804496290;
    11'd887: brom_out <= 64'd1153272281477598078;
    11'd247: brom_out <= 64'd3079117042164723820;
    11'd759: brom_out <= 64'd1885157749448756501;
    11'd503: brom_out <= 64'd287410934104796108;
    11'd1015: brom_out <= 64'd25262004549807233;
    11'd15: brom_out <= 64'd4373906864111961192;
    11'd527: brom_out <= 64'd5581925567248425011;
    11'd271: brom_out <= 64'd6143752504496732708;
    11'd783: brom_out <= 64'd8078411340332537200;
    11'd143: brom_out <= 64'd3405667996999341347;
    11'd655: brom_out <= 64'd8356640971005957295;
    11'd399: brom_out <= 64'd2937264643500724946;
    11'd911: brom_out <= 64'd7678224205154604892;
    11'd79: brom_out <= 64'd991733121096816246;
    11'd591: brom_out <= 64'd8206033862314336179;
    11'd335: brom_out <= 64'd5129160045159717183;
    11'd847: brom_out <= 64'd2359479212055339028;
    11'd207: brom_out <= 64'd964260620430079549;
    11'd719: brom_out <= 64'd281616783970276541;
    11'd463: brom_out <= 64'd7657127696980843717;
    11'd975: brom_out <= 64'd5088451844637495064;
    11'd47: brom_out <= 64'd1674291621165505607;
    11'd559: brom_out <= 64'd7402170804642201058;
    11'd303: brom_out <= 64'd3049253393215885299;
    11'd815: brom_out <= 64'd1572212746857595784;
    11'd175: brom_out <= 64'd4523172126112293441;
    11'd687: brom_out <= 64'd5471432485527519578;
    11'd431: brom_out <= 64'd968559680937005248;
    11'd943: brom_out <= 64'd8674281730199549271;
    11'd111: brom_out <= 64'd7186500760229875053;
    11'd623: brom_out <= 64'd7912654433847146065;
    11'd367: brom_out <= 64'd2944315729599332973;
    11'd879: brom_out <= 64'd6279407103230115525;
    11'd239: brom_out <= 64'd7701025136151381857;
    11'd751: brom_out <= 64'd3167893952487493944;
    11'd495: brom_out <= 64'd693939813520258859;
    11'd1007: brom_out <= 64'd8065342724630909459;
    11'd31: brom_out <= 64'd5596293620407173703;
    11'd543: brom_out <= 64'd5417023988817079832;
    11'd287: brom_out <= 64'd6615395692181224670;
    11'd799: brom_out <= 64'd8810587607558976549;
    11'd159: brom_out <= 64'd8308116381684268102;
    11'd671: brom_out <= 64'd4756412739101574244;
    11'd415: brom_out <= 64'd2099379525012808838;
    11'd927: brom_out <= 64'd3079009539254210979;
    11'd95: brom_out <= 64'd7138994063059429231;
    11'd607: brom_out <= 64'd7804553392680594608;
    11'd351: brom_out <= 64'd6867301955756113651;
    11'd863: brom_out <= 64'd3486478549657754942;
    11'd223: brom_out <= 64'd7442965855326153148;
    11'd735: brom_out <= 64'd3314498144052701739;
    11'd479: brom_out <= 64'd3294907764858559824;
    11'd991: brom_out <= 64'd315347814386475463;
    11'd63: brom_out <= 64'd8674474176990565409;
    11'd575: brom_out <= 64'd4463176173192127330;
    11'd319: brom_out <= 64'd5346911085079280798;
    11'd831: brom_out <= 64'd3850279675568096104;
    11'd191: brom_out <= 64'd1549853121982486025;
    11'd703: brom_out <= 64'd448403919027889030;
    11'd447: brom_out <= 64'd8460182789291736091;
    11'd959: brom_out <= 64'd1320547198527024793;
    11'd127: brom_out <= 64'd1680679157528580243;
    11'd639: brom_out <= 64'd5602381032211604622;
    11'd383: brom_out <= 64'd1405441374437402737;
    11'd895: brom_out <= 64'd7708772373098359625;
    11'd255: brom_out <= 64'd8632183450091772719;
    11'd767: brom_out <= 64'd6055970653617461320;
    11'd511: brom_out <= 64'd631785061731105457;
    11'd1023: brom_out <= 64'd9068072491154627648;
    default: brom_out <= 64'h1;
    endcase
end

generate
    if(DELAY == 1) begin
        assign b = brom_out;
    end
endgenerate

endmodule

//-------------------------------------------------------------------------------------------------

module tw_rom_11_ntt_nwc
#(
    parameter LOGN  = 11,
    parameter LOGQ  = 64,
    parameter DELAY = 1,
    parameter STAGE = 11
)(
    input            clk,
    input [LOGN-1:0] raddr,
    output[LOGQ-1:0] b
);

(* ram_style = "block" *)
reg [LOGQ-1:0] brom_out, brom_out2;

always @(posedge clk) begin
    case(raddr[STAGE-1:0])
    12'd0: brom_out <= 64'd3123572105583683402;
    12'd1024: brom_out <= 64'd6210072964040673020;
    12'd512: brom_out <= 64'd3342237017047793373;
    12'd1536: brom_out <= 64'd7355277617520634586;
    12'd256: brom_out <= 64'd3731688155441134519;
    12'd1280: brom_out <= 64'd746197257148082134;
    12'd768: brom_out <= 64'd6882017126725196445;
    12'd1792: brom_out <= 64'd2557864372178560436;
    12'd128: brom_out <= 64'd2166440950627386257;
    12'd1152: brom_out <= 64'd4591221540589937516;
    12'd640: brom_out <= 64'd7716981219181600943;
    12'd1664: brom_out <= 64'd2189049372073667650;
    12'd384: brom_out <= 64'd2311612871753849791;
    12'd1408: brom_out <= 64'd4072019081843533474;
    12'd896: brom_out <= 64'd8712181218839813404;
    12'd1920: brom_out <= 64'd6857881424320852643;
    12'd64: brom_out <= 64'd8494350379341673211;
    12'd1088: brom_out <= 64'd1450015595554632774;
    12'd576: brom_out <= 64'd7549463873573661007;
    12'd1600: brom_out <= 64'd1233914361232676098;
    12'd320: brom_out <= 64'd886198867756178430;
    12'd1344: brom_out <= 64'd1956066437631741368;
    12'd832: brom_out <= 64'd5627149728544187386;
    12'd1856: brom_out <= 64'd8274937244593370322;
    12'd192: brom_out <= 64'd7988979667361662759;
    12'd1216: brom_out <= 64'd4666592458098914089;
    12'd704: brom_out <= 64'd1298045902539398265;
    12'd1728: brom_out <= 64'd1761611861532361913;
    12'd448: brom_out <= 64'd5180878151982048690;
    12'd1472: brom_out <= 64'd4469892064000190110;
    12'd960: brom_out <= 64'd6523866588431288244;
    12'd1984: brom_out <= 64'd3574342989557969396;
    12'd32: brom_out <= 64'd2297192634176996362;
    12'd1056: brom_out <= 64'd6069782419959589417;
    12'd544: brom_out <= 64'd1646706165409496394;
    12'd1568: brom_out <= 64'd523334166551111434;
    12'd288: brom_out <= 64'd1919750695143281821;
    12'd1312: brom_out <= 64'd2442056004070379668;
    12'd800: brom_out <= 64'd750627169207456669;
    12'd1824: brom_out <= 64'd4993004925835321305;
    12'd160: brom_out <= 64'd2241191925486500147;
    12'd1184: brom_out <= 64'd458410435875458368;
    12'd672: brom_out <= 64'd8086341980048887515;
    12'd1696: brom_out <= 64'd6003204951930659681;
    12'd416: brom_out <= 64'd3385433203628413105;
    12'd1440: brom_out <= 64'd8492664244705889703;
    12'd928: brom_out <= 64'd4372975299754604474;
    12'd1952: brom_out <= 64'd6390291119259659044;
    12'd96: brom_out <= 64'd2044384050544942103;
    12'd1120: brom_out <= 64'd9137343943776462522;
    12'd608: brom_out <= 64'd8385457506386328156;
    12'd1632: brom_out <= 64'd7245898508682997123;
    12'd352: brom_out <= 64'd3936095812733887896;
    12'd1376: brom_out <= 64'd6175264778840526681;
    12'd864: brom_out <= 64'd6278320169781233282;
    12'd1888: brom_out <= 64'd1131343834085286502;
    12'd224: brom_out <= 64'd1067021338766054600;
    12'd1248: brom_out <= 64'd6708377314894467913;
    12'd736: brom_out <= 64'd448441719830181284;
    12'd1760: brom_out <= 64'd3462450930575773083;
    12'd480: brom_out <= 64'd2053072489035715110;
    12'd1504: brom_out <= 64'd3571446628147881729;
    12'd992: brom_out <= 64'd3266189979002004855;
    12'd2016: brom_out <= 64'd420841380367849997;
    12'd16: brom_out <= 64'd783182616177207598;
    12'd1040: brom_out <= 64'd2234302429879756578;
    12'd528: brom_out <= 64'd3991548750242451139;
    12'd1552: brom_out <= 64'd8692922177817170600;
    12'd272: brom_out <= 64'd1385594427132341856;
    12'd1296: brom_out <= 64'd8603143574189759185;
    12'd784: brom_out <= 64'd5359476522671379006;
    12'd1808: brom_out <= 64'd5881082224657863024;
    12'd144: brom_out <= 64'd8678182383998953170;
    12'd1168: brom_out <= 64'd3272127048956024083;
    12'd656: brom_out <= 64'd4701785531912350872;
    12'd1680: brom_out <= 64'd6626025465408209031;
    12'd400: brom_out <= 64'd3629578186473598833;
    12'd1424: brom_out <= 64'd3675762244302706408;
    12'd912: brom_out <= 64'd3735955948613914669;
    12'd1936: brom_out <= 64'd1957563335978200627;
    12'd80: brom_out <= 64'd4538474818802576657;
    12'd1104: brom_out <= 64'd6626597374803946101;
    12'd592: brom_out <= 64'd1697847849446268024;
    12'd1616: brom_out <= 64'd580163830187804849;
    12'd336: brom_out <= 64'd1568588832890587063;
    12'd1360: brom_out <= 64'd5321140009370534395;
    12'd848: brom_out <= 64'd909952118566978648;
    12'd1872: brom_out <= 64'd5254482570358799123;
    12'd208: brom_out <= 64'd2763390214731174683;
    12'd1232: brom_out <= 64'd833082138960878313;
    12'd720: brom_out <= 64'd6155954812303474773;
    12'd1744: brom_out <= 64'd2216879211519118055;
    12'd464: brom_out <= 64'd2896518042700706045;
    12'd1488: brom_out <= 64'd7856169405632948213;
    12'd976: brom_out <= 64'd5955208306166495403;
    12'd2000: brom_out <= 64'd2054155455637453233;
    12'd48: brom_out <= 64'd7090515701415971787;
    12'd1072: brom_out <= 64'd5471267595669168738;
    12'd560: brom_out <= 64'd2185353284342592968;
    12'd1584: brom_out <= 64'd7169004200705162714;
    12'd304: brom_out <= 64'd6956973355261008306;
    12'd1328: brom_out <= 64'd8302364376193292339;
    12'd816: brom_out <= 64'd286212631758874401;
    12'd1840: brom_out <= 64'd4906289506850021489;
    12'd176: brom_out <= 64'd1731669540915554494;
    12'd1200: brom_out <= 64'd7390300012921230879;
    12'd688: brom_out <= 64'd2343288219589085431;
    12'd1712: brom_out <= 64'd3124729955377220718;
    12'd432: brom_out <= 64'd339695076337037417;
    12'd1456: brom_out <= 64'd5872896871016669062;
    12'd944: brom_out <= 64'd7281917613505427323;
    12'd1968: brom_out <= 64'd1566986677748489042;
    12'd112: brom_out <= 64'd1942395595740367878;
    12'd1136: brom_out <= 64'd8781926067352473327;
    12'd624: brom_out <= 64'd2316648801153845325;
    12'd1648: brom_out <= 64'd8602699726710703741;
    12'd368: brom_out <= 64'd7791825354405238667;
    12'd1392: brom_out <= 64'd3439357931940964981;
    12'd880: brom_out <= 64'd726214298144433543;
    12'd1904: brom_out <= 64'd8061057984538643763;
    12'd240: brom_out <= 64'd3273602566738736569;
    12'd1264: brom_out <= 64'd7095699506140280224;
    12'd752: brom_out <= 64'd8893004132663739787;
    12'd1776: brom_out <= 64'd7930634006186368289;
    12'd496: brom_out <= 64'd4243592479602137596;
    12'd1520: brom_out <= 64'd8597286734662722249;
    12'd1008: brom_out <= 64'd6451814558501019995;
    12'd2032: brom_out <= 64'd9070399929026337210;
    12'd8: brom_out <= 64'd9116887236292092934;
    12'd1032: brom_out <= 64'd1606426951588592996;
    12'd520: brom_out <= 64'd4861487013059270599;
    12'd1544: brom_out <= 64'd260102973946485741;
    12'd264: brom_out <= 64'd5773698677946619728;
    12'd1288: brom_out <= 64'd4103816905759410609;
    12'd776: brom_out <= 64'd6892261297693813742;
    12'd1800: brom_out <= 64'd6333188063536259820;
    12'd136: brom_out <= 64'd7381661895931309007;
    12'd1160: brom_out <= 64'd5603901911539001522;
    12'd648: brom_out <= 64'd533005732002511292;
    12'd1672: brom_out <= 64'd7569204040891336436;
    12'd392: brom_out <= 64'd8057244330901810898;
    12'd1416: brom_out <= 64'd3214535847531560904;
    12'd904: brom_out <= 64'd4952848716949994613;
    12'd1928: brom_out <= 64'd6248621890190537167;
    12'd72: brom_out <= 64'd8874707211531011500;
    12'd1096: brom_out <= 64'd7427856066069298956;
    12'd584: brom_out <= 64'd603888116924036094;
    12'd1608: brom_out <= 64'd2754644077759772339;
    12'd328: brom_out <= 64'd9095063640756157767;
    12'd1352: brom_out <= 64'd632859793328261011;
    12'd840: brom_out <= 64'd6630697316414989991;
    12'd1864: brom_out <= 64'd3752299925704190949;
    12'd200: brom_out <= 64'd9198323919124624838;
    12'd1224: brom_out <= 64'd1874950184072912965;
    12'd712: brom_out <= 64'd2715642996503054597;
    12'd1736: brom_out <= 64'd308955336635552488;
    12'd456: brom_out <= 64'd2245186807235680102;
    12'd1480: brom_out <= 64'd4172640202111168758;
    12'd968: brom_out <= 64'd4077182461502919803;
    12'd1992: brom_out <= 64'd2732141223331029993;
    12'd40: brom_out <= 64'd2878487246493840219;
    12'd1064: brom_out <= 64'd660030551745809489;
    12'd552: brom_out <= 64'd3791309886402846957;
    12'd1576: brom_out <= 64'd1017928595862416507;
    12'd296: brom_out <= 64'd2442907485869086535;
    12'd1320: brom_out <= 64'd2849457659749957061;
    12'd808: brom_out <= 64'd7900749707574746965;
    12'd1832: brom_out <= 64'd8078662181464149966;
    12'd168: brom_out <= 64'd3176271261472844478;
    12'd1192: brom_out <= 64'd6464813145287066772;
    12'd680: brom_out <= 64'd950537228048801516;
    12'd1704: brom_out <= 64'd5831342265267309707;
    12'd424: brom_out <= 64'd4289164553228020220;
    12'd1448: brom_out <= 64'd5288258242696056923;
    12'd936: brom_out <= 64'd525250263869464149;
    12'd1960: brom_out <= 64'd7174949674258229829;
    12'd104: brom_out <= 64'd6622200784980244722;
    12'd1128: brom_out <= 64'd5197744071544625781;
    12'd616: brom_out <= 64'd1870963276953716576;
    12'd1640: brom_out <= 64'd895301291553104279;
    12'd360: brom_out <= 64'd3677393688610455850;
    12'd1384: brom_out <= 64'd3848288126021735160;
    12'd872: brom_out <= 64'd8876519078171770475;
    12'd1896: brom_out <= 64'd8501762627247681237;
    12'd232: brom_out <= 64'd3844352581851178287;
    12'd1256: brom_out <= 64'd375583526895939806;
    12'd744: brom_out <= 64'd4227784374869932528;
    12'd1768: brom_out <= 64'd3055783759957392061;
    12'd488: brom_out <= 64'd2128126771058898294;
    12'd1512: brom_out <= 64'd8955842841681352102;
    12'd1000: brom_out <= 64'd5723458789648090611;
    12'd2024: brom_out <= 64'd2741046798909788638;
    12'd24: brom_out <= 64'd344236587637152853;
    12'd1048: brom_out <= 64'd2942695266708798427;
    12'd536: brom_out <= 64'd7569686600946786322;
    12'd1560: brom_out <= 64'd1387079546863439318;
    12'd280: brom_out <= 64'd8883051673035921128;
    12'd1304: brom_out <= 64'd3306537775828484712;
    12'd792: brom_out <= 64'd6277976730879919786;
    12'd1816: brom_out <= 64'd7623086500210741289;
    12'd152: brom_out <= 64'd9176452086153447835;
    12'd1176: brom_out <= 64'd918690905556436854;
    12'd664: brom_out <= 64'd5533029577537463138;
    12'd1688: brom_out <= 64'd4203409571678735110;
    12'd408: brom_out <= 64'd1933131145020944084;
    12'd1432: brom_out <= 64'd949940012474322966;
    12'd920: brom_out <= 64'd2805883654978644739;
    12'd1944: brom_out <= 64'd5706782360995185956;
    12'd88: brom_out <= 64'd3318477840404178090;
    12'd1112: brom_out <= 64'd7321808279184263451;
    12'd600: brom_out <= 64'd8092842424723859072;
    12'd1624: brom_out <= 64'd7632207296033674789;
    12'd344: brom_out <= 64'd7913275755520123680;
    12'd1368: brom_out <= 64'd405464615108494398;
    12'd856: brom_out <= 64'd2379697201198083169;
    12'd1880: brom_out <= 64'd3839550017271574187;
    12'd216: brom_out <= 64'd3761537950009634296;
    12'd1240: brom_out <= 64'd5373508937008256770;
    12'd728: brom_out <= 64'd5367381007592077200;
    12'd1752: brom_out <= 64'd2818325502700138116;
    12'd472: brom_out <= 64'd583488639536759707;
    12'd1496: brom_out <= 64'd4265007619178284370;
    12'd984: brom_out <= 64'd7168872089427602820;
    12'd2008: brom_out <= 64'd345357047224859191;
    12'd56: brom_out <= 64'd1086385232282484544;
    12'd1080: brom_out <= 64'd7947286727604420409;
    12'd568: brom_out <= 64'd2330276115058745628;
    12'd1592: brom_out <= 64'd3736964995834394654;
    12'd312: brom_out <= 64'd2804869329954832515;
    12'd1336: brom_out <= 64'd7493287858764811070;
    12'd824: brom_out <= 64'd4900828823461895728;
    12'd1848: brom_out <= 64'd9098226647448061870;
    12'd184: brom_out <= 64'd6954178270385628264;
    12'd1208: brom_out <= 64'd4803907488525433514;
    12'd696: brom_out <= 64'd5307950595005733108;
    12'd1720: brom_out <= 64'd4480820987357422708;
    12'd440: brom_out <= 64'd3543156659599247151;
    12'd1464: brom_out <= 64'd1665907952920558564;
    12'd952: brom_out <= 64'd6982166819690192683;
    12'd1976: brom_out <= 64'd3434616805118562592;
    12'd120: brom_out <= 64'd1553290069140339772;
    12'd1144: brom_out <= 64'd490458484326936661;
    12'd632: brom_out <= 64'd2799746443987803563;
    12'd1656: brom_out <= 64'd950581874849829949;
    12'd376: brom_out <= 64'd7421368905880236143;
    12'd1400: brom_out <= 64'd141354680560203362;
    12'd888: brom_out <= 64'd761161538639400956;
    12'd1912: brom_out <= 64'd3771997065343949633;
    12'd248: brom_out <= 64'd4963424960183830701;
    12'd1272: brom_out <= 64'd5831912821561222187;
    12'd760: brom_out <= 64'd7821115560719082390;
    12'd1784: brom_out <= 64'd8463071353887895632;
    12'd504: brom_out <= 64'd1920259732134664347;
    12'd1528: brom_out <= 64'd6950438028055682140;
    12'd1016: brom_out <= 64'd6774251290066746706;
    12'd2040: brom_out <= 64'd1423492101511112774;
    12'd4: brom_out <= 64'd1594287808237617298;
    12'd1028: brom_out <= 64'd1950883529623070579;
    12'd516: brom_out <= 64'd8872362742624299435;
    12'd1540: brom_out <= 64'd6105195955178212147;
    12'd260: brom_out <= 64'd902376913565620621;
    12'd1284: brom_out <= 64'd2384214784490016440;
    12'd772: brom_out <= 64'd349749007813654970;
    12'd1796: brom_out <= 64'd8280723915928495026;
    12'd132: brom_out <= 64'd6006429786082668144;
    12'd1156: brom_out <= 64'd87775309465218771;
    12'd644: brom_out <= 64'd6507524922779195206;
    12'd1668: brom_out <= 64'd1170532761557822926;
    12'd388: brom_out <= 64'd9061822383527925634;
    12'd1412: brom_out <= 64'd5973400624239486279;
    12'd900: brom_out <= 64'd4956123448797288985;
    12'd1924: brom_out <= 64'd104829509605271681;
    12'd68: brom_out <= 64'd4447161808775547377;
    12'd1092: brom_out <= 64'd8263840048186713893;
    12'd580: brom_out <= 64'd3723614080956210237;
    12'd1604: brom_out <= 64'd2106133836070735714;
    12'd324: brom_out <= 64'd5954126167444784680;
    12'd1348: brom_out <= 64'd5837535850480979167;
    12'd836: brom_out <= 64'd2032034460964293559;
    12'd1860: brom_out <= 64'd6799933047304790248;
    12'd196: brom_out <= 64'd5944579320629495743;
    12'd1220: brom_out <= 64'd1114328369126443520;
    12'd708: brom_out <= 64'd3210665055033323269;
    12'd1732: brom_out <= 64'd331662582474243093;
    12'd452: brom_out <= 64'd7285995299631463365;
    12'd1476: brom_out <= 64'd5591146297170291876;
    12'd964: brom_out <= 64'd2927030839530446166;
    12'd1988: brom_out <= 64'd9180053981269946509;
    12'd36: brom_out <= 64'd2038400528523470856;
    12'd1060: brom_out <= 64'd4945910978679130052;
    12'd548: brom_out <= 64'd3322412654452468391;
    12'd1572: brom_out <= 64'd6955311913223503755;
    12'd292: brom_out <= 64'd6714396605823359954;
    12'd1316: brom_out <= 64'd6762723344434804777;
    12'd804: brom_out <= 64'd631431952861437530;
    12'd1828: brom_out <= 64'd6502067971870131402;
    12'd164: brom_out <= 64'd7056313233161554884;
    12'd1188: brom_out <= 64'd5508599142792187880;
    12'd676: brom_out <= 64'd8117785985794032769;
    12'd1700: brom_out <= 64'd7189340714624472391;
    12'd420: brom_out <= 64'd8077247110993010098;
    12'd1444: brom_out <= 64'd385434811086117404;
    12'd932: brom_out <= 64'd6140272816859085023;
    12'd1956: brom_out <= 64'd4093413828459857685;
    12'd100: brom_out <= 64'd7212496672846126617;
    12'd1124: brom_out <= 64'd4716495894692356985;
    12'd612: brom_out <= 64'd8861948288597181352;
    12'd1636: brom_out <= 64'd7997500746202064856;
    12'd356: brom_out <= 64'd7036761341881640631;
    12'd1380: brom_out <= 64'd373931093920173974;
    12'd868: brom_out <= 64'd8672482648636030314;
    12'd1892: brom_out <= 64'd2735304322641470733;
    12'd228: brom_out <= 64'd8322563467653039148;
    12'd1252: brom_out <= 64'd5402537941179410779;
    12'd740: brom_out <= 64'd7443079129547343031;
    12'd1764: brom_out <= 64'd9213216472849345386;
    12'd484: brom_out <= 64'd4256246873122223388;
    12'd1508: brom_out <= 64'd4867178542899370437;
    12'd996: brom_out <= 64'd2117247787424601565;
    12'd2020: brom_out <= 64'd8548194336979807;
    12'd20: brom_out <= 64'd84178952316759680;
    12'd1044: brom_out <= 64'd8460257235923533062;
    12'd532: brom_out <= 64'd5332876089822586158;
    12'd1556: brom_out <= 64'd8505599904453139329;
    12'd276: brom_out <= 64'd3777627475796403316;
    12'd1300: brom_out <= 64'd6674428628901193372;
    12'd788: brom_out <= 64'd500810411488742958;
    12'd1812: brom_out <= 64'd7041229430920456324;
    12'd148: brom_out <= 64'd412180794031832049;
    12'd1172: brom_out <= 64'd7597615280424166823;
    12'd660: brom_out <= 64'd7986399044849774194;
    12'd1684: brom_out <= 64'd8682695751401982685;
    12'd404: brom_out <= 64'd361526547022696037;
    12'd1428: brom_out <= 64'd4511931667639884277;
    12'd916: brom_out <= 64'd6418507330796271220;
    12'd1940: brom_out <= 64'd6263587321880250693;
    12'd84: brom_out <= 64'd4993034077449917730;
    12'd1108: brom_out <= 64'd589228948138830458;
    12'd596: brom_out <= 64'd8434086446192677801;
    12'd1620: brom_out <= 64'd3496472476864176797;
    12'd340: brom_out <= 64'd5182291076888013309;
    12'd1364: brom_out <= 64'd3505693018995845744;
    12'd852: brom_out <= 64'd647644701333757196;
    12'd1876: brom_out <= 64'd9115268039952312342;
    12'd212: brom_out <= 64'd6713049577875831491;
    12'd1236: brom_out <= 64'd6078949513059548796;
    12'd724: brom_out <= 64'd8731838398833267099;
    12'd1748: brom_out <= 64'd381924365733082925;
    12'd468: brom_out <= 64'd526278107207560948;
    12'd1492: brom_out <= 64'd6012936457007095415;
    12'd980: brom_out <= 64'd6179895911262856559;
    12'd2004: brom_out <= 64'd7105295964005438960;
    12'd52: brom_out <= 64'd5519475337282045668;
    12'd1076: brom_out <= 64'd5607239368114546459;
    12'd564: brom_out <= 64'd8137793089463064705;
    12'd1588: brom_out <= 64'd2621261092389224257;
    12'd308: brom_out <= 64'd140754322501936048;
    12'd1332: brom_out <= 64'd2731388838744875166;
    12'd820: brom_out <= 64'd5500938849019406519;
    12'd1844: brom_out <= 64'd9002304854898473773;
    12'd180: brom_out <= 64'd8488516030236336871;
    12'd1204: brom_out <= 64'd1581299506068635164;
    12'd692: brom_out <= 64'd8426404365643318269;
    12'd1716: brom_out <= 64'd6086578453601839060;
    12'd436: brom_out <= 64'd3958099533337224045;
    12'd1460: brom_out <= 64'd7981229849417595750;
    12'd948: brom_out <= 64'd6960988389091375728;
    12'd1972: brom_out <= 64'd4665671487038613092;
    12'd116: brom_out <= 64'd2682137270946396050;
    12'd1140: brom_out <= 64'd447817529184977423;
    12'd628: brom_out <= 64'd367318817448002619;
    12'd1652: brom_out <= 64'd1051387047755393606;
    12'd372: brom_out <= 64'd1691932192495541122;
    12'd1396: brom_out <= 64'd957899819091921531;
    12'd884: brom_out <= 64'd1524891256519788450;
    12'd1908: brom_out <= 64'd5505288545782259845;
    12'd244: brom_out <= 64'd7379185160575291364;
    12'd1268: brom_out <= 64'd3878416946790585359;
    12'd756: brom_out <= 64'd3824227222565397005;
    12'd1780: brom_out <= 64'd6444946389109126637;
    12'd500: brom_out <= 64'd3487447292574180815;
    12'd1524: brom_out <= 64'd1918271444866228967;
    12'd1012: brom_out <= 64'd7031234002988880400;
    12'd2036: brom_out <= 64'd2112615497361464837;
    12'd12: brom_out <= 64'd2795111693195155866;
    12'd1036: brom_out <= 64'd472421530302321434;
    12'd524: brom_out <= 64'd6068520444408022295;
    12'd1548: brom_out <= 64'd1617224231272278262;
    12'd268: brom_out <= 64'd2569904008316410260;
    12'd1292: brom_out <= 64'd8526219922781128460;
    12'd780: brom_out <= 64'd8327465683114700851;
    12'd1804: brom_out <= 64'd7568443072540426724;
    12'd140: brom_out <= 64'd4629020314711264699;
    12'd1164: brom_out <= 64'd4332603151624655979;
    12'd652: brom_out <= 64'd3127355264627254150;
    12'd1676: brom_out <= 64'd9033233996773343847;
    12'd396: brom_out <= 64'd9005688290792999644;
    12'd1420: brom_out <= 64'd6030955605040008120;
    12'd908: brom_out <= 64'd8789643826458638393;
    12'd1932: brom_out <= 64'd7552849624034460758;
    12'd76: brom_out <= 64'd6162735083455312198;
    12'd1100: brom_out <= 64'd6524744156397851803;
    12'd588: brom_out <= 64'd5579413719146707083;
    12'd1612: brom_out <= 64'd948297851783343744;
    12'd332: brom_out <= 64'd81185299302372879;
    12'd1356: brom_out <= 64'd3063166609615503984;
    12'd844: brom_out <= 64'd795649999775240663;
    12'd1868: brom_out <= 64'd8037251786593648802;
    12'd204: brom_out <= 64'd502777772910858913;
    12'd1228: brom_out <= 64'd6597444450441397719;
    12'd716: brom_out <= 64'd5846223268732879046;
    12'd1740: brom_out <= 64'd6130050090479151203;
    12'd460: brom_out <= 64'd2384975474288463368;
    12'd1484: brom_out <= 64'd3596112534661279898;
    12'd972: brom_out <= 64'd7221494124396180503;
    12'd1996: brom_out <= 64'd4605276482808534409;
    12'd44: brom_out <= 64'd2944422568018111881;
    12'd1068: brom_out <= 64'd3605998430247226191;
    12'd556: brom_out <= 64'd1587569415606107148;
    12'd1580: brom_out <= 64'd760642633244382233;
    12'd300: brom_out <= 64'd4815585788747747930;
    12'd1324: brom_out <= 64'd4659110683430105708;
    12'd812: brom_out <= 64'd7686812788309527859;
    12'd1836: brom_out <= 64'd3110662909970991713;
    12'd172: brom_out <= 64'd7674152101976600121;
    12'd1196: brom_out <= 64'd4635868544219197072;
    12'd684: brom_out <= 64'd4116964532439010750;
    12'd1708: brom_out <= 64'd5080690067356352286;
    12'd428: brom_out <= 64'd3101728032514437051;
    12'd1452: brom_out <= 64'd8115736187040631118;
    12'd940: brom_out <= 64'd8187738356454920847;
    12'd1964: brom_out <= 64'd5730693877087875771;
    12'd108: brom_out <= 64'd5610169279134306168;
    12'd1132: brom_out <= 64'd4612706075332010148;
    12'd620: brom_out <= 64'd3229527714353233405;
    12'd1644: brom_out <= 64'd6366856511970655221;
    12'd364: brom_out <= 64'd9028424703745913643;
    12'd1388: brom_out <= 64'd2612253775413894197;
    12'd876: brom_out <= 64'd9058913656626322415;
    12'd1900: brom_out <= 64'd5884626759484195837;
    12'd236: brom_out <= 64'd1976917306024987061;
    12'd1260: brom_out <= 64'd3928066874472912805;
    12'd748: brom_out <= 64'd8249885220722612302;
    12'd1772: brom_out <= 64'd3528258301290806711;
    12'd492: brom_out <= 64'd1657488472428570923;
    12'd1516: brom_out <= 64'd3821666041687242524;
    12'd1004: brom_out <= 64'd6416282645049431358;
    12'd2028: brom_out <= 64'd4862535682100292549;
    12'd28: brom_out <= 64'd5409368920540923008;
    12'd1052: brom_out <= 64'd4009441914452456916;
    12'd540: brom_out <= 64'd3408413532395370996;
    12'd1564: brom_out <= 64'd8028084994748216739;
    12'd284: brom_out <= 64'd3849333415702798784;
    12'd1308: brom_out <= 64'd8365722423632335032;
    12'd796: brom_out <= 64'd3427611725193605315;
    12'd1820: brom_out <= 64'd7864825205091798631;
    12'd156: brom_out <= 64'd5396538137592370747;
    12'd1180: brom_out <= 64'd43072760317062206;
    12'd668: brom_out <= 64'd2982463332641780795;
    12'd1692: brom_out <= 64'd2491406867419859581;
    12'd412: brom_out <= 64'd4447550820321395770;
    12'd1436: brom_out <= 64'd5801594966488479138;
    12'd924: brom_out <= 64'd7852199942964421451;
    12'd1948: brom_out <= 64'd4178440991420012237;
    12'd92: brom_out <= 64'd6952270401479331297;
    12'd1116: brom_out <= 64'd4578300779314317085;
    12'd604: brom_out <= 64'd924172865789957521;
    12'd1628: brom_out <= 64'd5688887396703162594;
    12'd348: brom_out <= 64'd2748649208425336417;
    12'd1372: brom_out <= 64'd7049664898306437476;
    12'd860: brom_out <= 64'd4747326262452797291;
    12'd1884: brom_out <= 64'd985147216069003303;
    12'd220: brom_out <= 64'd4813892700286973804;
    12'd1244: brom_out <= 64'd1259792959611445980;
    12'd732: brom_out <= 64'd6053220151492819634;
    12'd1756: brom_out <= 64'd8508099142022419643;
    12'd476: brom_out <= 64'd8371120847098266361;
    12'd1500: brom_out <= 64'd7772347693311743621;
    12'd988: brom_out <= 64'd563604324382919887;
    12'd2012: brom_out <= 64'd5439372450993987387;
    12'd60: brom_out <= 64'd231306203269935887;
    12'd1084: brom_out <= 64'd6612377017870351741;
    12'd572: brom_out <= 64'd3388949387369608667;
    12'd1596: brom_out <= 64'd8106844442911889453;
    12'd316: brom_out <= 64'd777497982063491819;
    12'd1340: brom_out <= 64'd8985719704801141523;
    12'd828: brom_out <= 64'd1555620882056217295;
    12'd1852: brom_out <= 64'd2881664385376323498;
    12'd188: brom_out <= 64'd3336878337925885369;
    12'd1212: brom_out <= 64'd1009851933266404927;
    12'd700: brom_out <= 64'd9202131982711188586;
    12'd1724: brom_out <= 64'd3231135258943435442;
    12'd444: brom_out <= 64'd4061131916105246763;
    12'd1468: brom_out <= 64'd5593127481509872288;
    12'd956: brom_out <= 64'd5215064358567618019;
    12'd1980: brom_out <= 64'd4564263216878088566;
    12'd124: brom_out <= 64'd8265708178362476224;
    12'd1148: brom_out <= 64'd6596969282323087897;
    12'd636: brom_out <= 64'd4294714109527455000;
    12'd1660: brom_out <= 64'd2395015109056088141;
    12'd380: brom_out <= 64'd403207746426225723;
    12'd1404: brom_out <= 64'd4069951574478518978;
    12'd892: brom_out <= 64'd4651171245899521217;
    12'd1916: brom_out <= 64'd6459172628559921705;
    12'd252: brom_out <= 64'd1146151887566287582;
    12'd1276: brom_out <= 64'd8859555029944229464;
    12'd764: brom_out <= 64'd7053943251416293791;
    12'd1788: brom_out <= 64'd92400884003435777;
    12'd508: brom_out <= 64'd3101654541177146791;
    12'd1532: brom_out <= 64'd6424226835471038558;
    12'd1020: brom_out <= 64'd5911746077465107851;
    12'd2044: brom_out <= 64'd3605580692623497747;
    12'd2: brom_out <= 64'd4161382131132605360;
    12'd1026: brom_out <= 64'd8294400354274293827;
    12'd514: brom_out <= 64'd4245248340976967157;
    12'd1538: brom_out <= 64'd7005760798045576267;
    12'd258: brom_out <= 64'd3125413967307849523;
    12'd1282: brom_out <= 64'd1354982801898793653;
    12'd770: brom_out <= 64'd5593298290473968207;
    12'd1794: brom_out <= 64'd7739085512538120589;
    12'd130: brom_out <= 64'd6427417093273440184;
    12'd1154: brom_out <= 64'd3808131466260275888;
    12'd642: brom_out <= 64'd1266239233228019763;
    12'd1666: brom_out <= 64'd7052090867174173971;
    12'd386: brom_out <= 64'd3616056455335921290;
    12'd1410: brom_out <= 64'd3148043341039269482;
    12'd898: brom_out <= 64'd2346589270844952759;
    12'd1922: brom_out <= 64'd6063326813558607448;
    12'd66: brom_out <= 64'd8735870872178958038;
    12'd1090: brom_out <= 64'd8799477870518799650;
    12'd578: brom_out <= 64'd5812217558536995975;
    12'd1602: brom_out <= 64'd7871887319621567624;
    12'd322: brom_out <= 64'd42305848928908451;
    12'd1346: brom_out <= 64'd513856896927873735;
    12'd834: brom_out <= 64'd1472777169665991434;
    12'd1858: brom_out <= 64'd2640221677355103899;
    12'd194: brom_out <= 64'd5166371174271619888;
    12'd1218: brom_out <= 64'd8433763352154848682;
    12'd706: brom_out <= 64'd5187949924568406697;
    12'd1730: brom_out <= 64'd6370911676719588588;
    12'd450: brom_out <= 64'd4030172962426199408;
    12'd1474: brom_out <= 64'd6778376992396069474;
    12'd962: brom_out <= 64'd1591397077274221089;
    12'd1986: brom_out <= 64'd7162683964198145608;
    12'd34: brom_out <= 64'd2539262627007689965;
    12'd1058: brom_out <= 64'd336401549822729772;
    12'd546: brom_out <= 64'd5998172594559044492;
    12'd1570: brom_out <= 64'd6478334644154555715;
    12'd290: brom_out <= 64'd6432916138033825836;
    12'd1314: brom_out <= 64'd2501962074965142941;
    12'd802: brom_out <= 64'd2317435503726077713;
    12'd1826: brom_out <= 64'd5235992488295912615;
    12'd162: brom_out <= 64'd7018917583447423622;
    12'd1186: brom_out <= 64'd3888056778530587651;
    12'd674: brom_out <= 64'd1708102970485337530;
    12'd1698: brom_out <= 64'd2851469000801802053;
    12'd418: brom_out <= 64'd7853994117985328905;
    12'd1442: brom_out <= 64'd3401575306703463020;
    12'd930: brom_out <= 64'd6877317548467700668;
    12'd1954: brom_out <= 64'd7103185062750783314;
    12'd98: brom_out <= 64'd5033644458990983072;
    12'd1122: brom_out <= 64'd4457221733501494314;
    12'd610: brom_out <= 64'd6901871725493421902;
    12'd1634: brom_out <= 64'd5811539893595560331;
    12'd354: brom_out <= 64'd3636856344111207334;
    12'd1378: brom_out <= 64'd5049677082286780231;
    12'd866: brom_out <= 64'd1256517597608267931;
    12'd1890: brom_out <= 64'd5807673899962685070;
    12'd226: brom_out <= 64'd3812088677365165897;
    12'd1250: brom_out <= 64'd8869517514595545325;
    12'd738: brom_out <= 64'd4547272604806793912;
    12'd1762: brom_out <= 64'd6121711115027851334;
    12'd482: brom_out <= 64'd869623750016964361;
    12'd1506: brom_out <= 64'd7538895155878924298;
    12'd994: brom_out <= 64'd2398707703947764450;
    12'd2018: brom_out <= 64'd3139470700951704937;
    12'd18: brom_out <= 64'd5291791690895949625;
    12'd1042: brom_out <= 64'd5504964789253506993;
    12'd530: brom_out <= 64'd2179428562918306485;
    12'd1554: brom_out <= 64'd3013380075501454019;
    12'd274: brom_out <= 64'd8320828789819456468;
    12'd1298: brom_out <= 64'd1244950926757250904;
    12'd786: brom_out <= 64'd177066268119183448;
    12'd1810: brom_out <= 64'd5754503534626256193;
    12'd146: brom_out <= 64'd6463543092520081206;
    12'd1170: brom_out <= 64'd7614153997158589913;
    12'd658: brom_out <= 64'd8427105068273902421;
    12'd1682: brom_out <= 64'd8763555563296182556;
    12'd402: brom_out <= 64'd6127895378780629091;
    12'd1426: brom_out <= 64'd6928605446208831427;
    12'd914: brom_out <= 64'd787612018681613361;
    12'd1938: brom_out <= 64'd7855429259490051967;
    12'd82: brom_out <= 64'd2219578339043977142;
    12'd1106: brom_out <= 64'd8713121753568537292;
    12'd594: brom_out <= 64'd8066481711723959380;
    12'd1618: brom_out <= 64'd7407469317649966302;
    12'd338: brom_out <= 64'd36977916334723084;
    12'd1362: brom_out <= 64'd7782935284441959380;
    12'd850: brom_out <= 64'd3602236584122824560;
    12'd1874: brom_out <= 64'd1021123098135788205;
    12'd210: brom_out <= 64'd8520131378825116961;
    12'd1234: brom_out <= 64'd1316765805752574193;
    12'd722: brom_out <= 64'd3205392293724576591;
    12'd1746: brom_out <= 64'd1143628808215917235;
    12'd466: brom_out <= 64'd8991850183852190750;
    12'd1490: brom_out <= 64'd9091022804974507130;
    12'd978: brom_out <= 64'd3088053723604747001;
    12'd2002: brom_out <= 64'd5623148121671206125;
    12'd50: brom_out <= 64'd7657043159525780525;
    12'd1074: brom_out <= 64'd8495822332160611203;
    12'd562: brom_out <= 64'd1679130689109720777;
    12'd1586: brom_out <= 64'd1568151740605117802;
    12'd306: brom_out <= 64'd3572451211808755669;
    12'd1330: brom_out <= 64'd3016753087757996057;
    12'd818: brom_out <= 64'd7409637591157424255;
    12'd1842: brom_out <= 64'd1327915948460867785;
    12'd178: brom_out <= 64'd5842552477701386526;
    12'd1202: brom_out <= 64'd4496194611457518364;
    12'd690: brom_out <= 64'd7462704917437603606;
    12'd1714: brom_out <= 64'd6366777947683303534;
    12'd434: brom_out <= 64'd6120561367020358740;
    12'd1458: brom_out <= 64'd6621892503978496011;
    12'd946: brom_out <= 64'd9046550912136285240;
    12'd1970: brom_out <= 64'd7201884348327293194;
    12'd114: brom_out <= 64'd767133063771333272;
    12'd1138: brom_out <= 64'd2561818334564375246;
    12'd626: brom_out <= 64'd5457559586433941288;
    12'd1650: brom_out <= 64'd1128788383963247148;
    12'd370: brom_out <= 64'd6413883711658996975;
    12'd1394: brom_out <= 64'd927205808884007408;
    12'd882: brom_out <= 64'd2283814024811077477;
    12'd1906: brom_out <= 64'd1342238341057611796;
    12'd242: brom_out <= 64'd6636571708981876228;
    12'd1266: brom_out <= 64'd5662731900612283352;
    12'd754: brom_out <= 64'd2567562405985803722;
    12'd1778: brom_out <= 64'd4735863391036245873;
    12'd498: brom_out <= 64'd3884633026447537169;
    12'd1522: brom_out <= 64'd2355835589563975467;
    12'd1010: brom_out <= 64'd8373242971525403027;
    12'd2034: brom_out <= 64'd8269699888498060215;
    12'd10: brom_out <= 64'd4607407384118149230;
    12'd1034: brom_out <= 64'd2782325799324638689;
    12'd522: brom_out <= 64'd5339941612673657853;
    12'd1546: brom_out <= 64'd2201871850899339104;
    12'd266: brom_out <= 64'd3709428719556243465;
    12'd1290: brom_out <= 64'd1585353406432777339;
    12'd778: brom_out <= 64'd4844702021110767552;
    12'd1802: brom_out <= 64'd1466922448770939007;
    12'd138: brom_out <= 64'd8263663049475472786;
    12'd1162: brom_out <= 64'd2437472423545569288;
    12'd650: brom_out <= 64'd1779378143287967658;
    12'd1674: brom_out <= 64'd5724966495240726420;
    12'd394: brom_out <= 64'd5773071269164981114;
    12'd1418: brom_out <= 64'd5932590464980392607;
    12'd906: brom_out <= 64'd7168388657041672505;
    12'd1930: brom_out <= 64'd381062116641522675;
    12'd74: brom_out <= 64'd811765929269079575;
    12'd1098: brom_out <= 64'd3784172596301817125;
    12'd586: brom_out <= 64'd3342083064961576527;
    12'd1610: brom_out <= 64'd2114146786529872706;
    12'd330: brom_out <= 64'd2580934252726307195;
    12'd1354: brom_out <= 64'd4059066379504251084;
    12'd842: brom_out <= 64'd6641457222189368918;
    12'd1866: brom_out <= 64'd8863909611002520133;
    12'd202: brom_out <= 64'd3079087207722465675;
    12'd1226: brom_out <= 64'd2827295680149049363;
    12'd714: brom_out <= 64'd5128305230030333456;
    12'd1738: brom_out <= 64'd5481820251577889089;
    12'd458: brom_out <= 64'd6307758981226501337;
    12'd1482: brom_out <= 64'd5812845803670824712;
    12'd970: brom_out <= 64'd4783216896920612281;
    12'd1994: brom_out <= 64'd5267121197034638085;
    12'd42: brom_out <= 64'd1841890384989310399;
    12'd1066: brom_out <= 64'd831002150678604344;
    12'd554: brom_out <= 64'd3069375341129563391;
    12'd1578: brom_out <= 64'd4344767874481239703;
    12'd298: brom_out <= 64'd7992055436492775547;
    12'd1322: brom_out <= 64'd6416667228388435455;
    12'd810: brom_out <= 64'd3091207899330601804;
    12'd1834: brom_out <= 64'd6627033872986159219;
    12'd170: brom_out <= 64'd6932390504227637120;
    12'd1194: brom_out <= 64'd2443508318932193909;
    12'd682: brom_out <= 64'd6081479337248015055;
    12'd1706: brom_out <= 64'd7764130815122539721;
    12'd426: brom_out <= 64'd6280175778077984849;
    12'd1450: brom_out <= 64'd6599130383498806289;
    12'd938: brom_out <= 64'd1252309368676415478;
    12'd1962: brom_out <= 64'd4480395508255192801;
    12'd106: brom_out <= 64'd3942996461323465180;
    12'd1130: brom_out <= 64'd4401921130714756231;
    12'd618: brom_out <= 64'd555821410683758034;
    12'd1642: brom_out <= 64'd5023515734586300393;
    12'd362: brom_out <= 64'd5526953088984257734;
    12'd1386: brom_out <= 64'd7815017051210755800;
    12'd874: brom_out <= 64'd1890273632003078815;
    12'd1898: brom_out <= 64'd5779175783193383990;
    12'd234: brom_out <= 64'd1456674837575388517;
    12'd1258: brom_out <= 64'd1418956800510201025;
    12'd746: brom_out <= 64'd7064874188067316261;
    12'd1770: brom_out <= 64'd1449330551565739163;
    12'd490: brom_out <= 64'd3215301725679354417;
    12'd1514: brom_out <= 64'd6558956959724034571;
    12'd1002: brom_out <= 64'd2930000210000861422;
    12'd2026: brom_out <= 64'd1463275534110631389;
    12'd26: brom_out <= 64'd1196098718942254763;
    12'd1050: brom_out <= 64'd8366114043396594506;
    12'd538: brom_out <= 64'd5984103877935957177;
    12'd1562: brom_out <= 64'd2949102692196058895;
    12'd282: brom_out <= 64'd7547575482964536409;
    12'd1306: brom_out <= 64'd3149938985678811660;
    12'd794: brom_out <= 64'd2002443587523568133;
    12'd1818: brom_out <= 64'd6668743251079113996;
    12'd154: brom_out <= 64'd5796109678201625407;
    12'd1178: brom_out <= 64'd1595342553448744058;
    12'd666: brom_out <= 64'd3519590871235660295;
    12'd1690: brom_out <= 64'd7458906364176709762;
    12'd410: brom_out <= 64'd8878971298747704074;
    12'd1434: brom_out <= 64'd3396121475613569590;
    12'd922: brom_out <= 64'd7365127815719282940;
    12'd1946: brom_out <= 64'd7606956865799178146;
    12'd90: brom_out <= 64'd2400666355134559122;
    12'd1114: brom_out <= 64'd8010437356180367926;
    12'd602: brom_out <= 64'd8758609324438474644;
    12'd1626: brom_out <= 64'd1146517788248817457;
    12'd346: brom_out <= 64'd3639190735179687537;
    12'd1370: brom_out <= 64'd5707924727106845397;
    12'd858: brom_out <= 64'd716495466631501188;
    12'd1882: brom_out <= 64'd6414603494018560970;
    12'd218: brom_out <= 64'd1592871631962342491;
    12'd1242: brom_out <= 64'd181668506279055852;
    12'd730: brom_out <= 64'd6744894345592053761;
    12'd1754: brom_out <= 64'd4037674446693902019;
    12'd474: brom_out <= 64'd5411874943025385150;
    12'd1498: brom_out <= 64'd359719403014682205;
    12'd986: brom_out <= 64'd24859528214763344;
    12'd2010: brom_out <= 64'd8119561780682838824;
    12'd58: brom_out <= 64'd6135325541824978667;
    12'd1082: brom_out <= 64'd4797535891935457436;
    12'd570: brom_out <= 64'd7241464595079900974;
    12'd1594: brom_out <= 64'd3606929189234260139;
    12'd314: brom_out <= 64'd7013113869652190949;
    12'd1338: brom_out <= 64'd1000493227257847315;
    12'd826: brom_out <= 64'd5333207141477065766;
    12'd1850: brom_out <= 64'd2869042744839996736;
    12'd186: brom_out <= 64'd8892600644819782934;
    12'd1210: brom_out <= 64'd1761679396632364677;
    12'd698: brom_out <= 64'd7486651560101348658;
    12'd1722: brom_out <= 64'd7901294082693364184;
    12'd442: brom_out <= 64'd1373994615435235519;
    12'd1466: brom_out <= 64'd6227174019170902624;
    12'd954: brom_out <= 64'd8831142828453098264;
    12'd1978: brom_out <= 64'd625727918417707050;
    12'd122: brom_out <= 64'd935707005244710622;
    12'd1146: brom_out <= 64'd1877248393457524943;
    12'd634: brom_out <= 64'd1316579341960321860;
    12'd1658: brom_out <= 64'd4191416174392406972;
    12'd378: brom_out <= 64'd8213979470788678857;
    12'd1402: brom_out <= 64'd4776594591265232375;
    12'd890: brom_out <= 64'd7289274910654307939;
    12'd1914: brom_out <= 64'd7098596105988351439;
    12'd250: brom_out <= 64'd8636431542623556342;
    12'd1274: brom_out <= 64'd2856467410577393100;
    12'd762: brom_out <= 64'd9057087941673552377;
    12'd1786: brom_out <= 64'd4724055599125808147;
    12'd506: brom_out <= 64'd7890148038881897550;
    12'd1530: brom_out <= 64'd4344459685671561063;
    12'd1018: brom_out <= 64'd1667366953149435079;
    12'd2042: brom_out <= 64'd5379642131606208872;
    12'd6: brom_out <= 64'd833853371947711770;
    12'd1030: brom_out <= 64'd889947342877147235;
    12'd518: brom_out <= 64'd3796405865253091106;
    12'd1542: brom_out <= 64'd6014537814613808573;
    12'd262: brom_out <= 64'd3826836417145052821;
    12'd1286: brom_out <= 64'd7609378528917516818;
    12'd774: brom_out <= 64'd9026635029389000381;
    12'd1798: brom_out <= 64'd8513140117475607861;
    12'd134: brom_out <= 64'd2192981460894983780;
    12'd1158: brom_out <= 64'd2717284282999342539;
    12'd646: brom_out <= 64'd5542434471175813321;
    12'd1670: brom_out <= 64'd2932745904589837228;
    12'd390: brom_out <= 64'd1077638811771035248;
    12'd1414: brom_out <= 64'd5547009549118445021;
    12'd902: brom_out <= 64'd3466959967303810227;
    12'd1926: brom_out <= 64'd1200663969910512904;
    12'd70: brom_out <= 64'd2930272707943786556;
    12'd1094: brom_out <= 64'd8535100517885305196;
    12'd582: brom_out <= 64'd2179382374964276344;
    12'd1606: brom_out <= 64'd7959052490157018496;
    12'd326: brom_out <= 64'd7160917862990901367;
    12'd1350: brom_out <= 64'd4870496060242192381;
    12'd838: brom_out <= 64'd2636451624071188702;
    12'd1862: brom_out <= 64'd517091244716182147;
    12'd198: brom_out <= 64'd8622631016638827589;
    12'd1222: brom_out <= 64'd7347896371767391775;
    12'd710: brom_out <= 64'd3178574472699619460;
    12'd1734: brom_out <= 64'd8901832433890731733;
    12'd454: brom_out <= 64'd2508667236487445379;
    12'd1478: brom_out <= 64'd2170222475619826595;
    12'd966: brom_out <= 64'd1812309815745216366;
    12'd1990: brom_out <= 64'd8692059923454255042;
    12'd38: brom_out <= 64'd6005123582676054331;
    12'd1062: brom_out <= 64'd255745229776933456;
    12'd550: brom_out <= 64'd71801563849700887;
    12'd1574: brom_out <= 64'd9044180726951058564;
    12'd294: brom_out <= 64'd5787202332160718093;
    12'd1318: brom_out <= 64'd5631415570082035830;
    12'd806: brom_out <= 64'd1590129923100941094;
    12'd1830: brom_out <= 64'd8418009426952650638;
    12'd166: brom_out <= 64'd6887211691168918066;
    12'd1190: brom_out <= 64'd3402428439857658913;
    12'd678: brom_out <= 64'd4359598444987897660;
    12'd1702: brom_out <= 64'd190397694499685176;
    12'd422: brom_out <= 64'd58494804674635643;
    12'd1446: brom_out <= 64'd9009490652745159817;
    12'd934: brom_out <= 64'd6766756384274140931;
    12'd1958: brom_out <= 64'd4599090932582395178;
    12'd102: brom_out <= 64'd9184521068795560933;
    12'd1126: brom_out <= 64'd6019436832580782773;
    12'd614: brom_out <= 64'd4424064624941582579;
    12'd1638: brom_out <= 64'd146279101367442789;
    12'd358: brom_out <= 64'd6313145164733755544;
    12'd1382: brom_out <= 64'd6833914128980402973;
    12'd870: brom_out <= 64'd3356671144027189909;
    12'd1894: brom_out <= 64'd1790287456568310240;
    12'd230: brom_out <= 64'd4624760394558543392;
    12'd1254: brom_out <= 64'd4305286141946115626;
    12'd742: brom_out <= 64'd8755047956121748583;
    12'd1766: brom_out <= 64'd162010141640127860;
    12'd486: brom_out <= 64'd2515444599521314796;
    12'd1510: brom_out <= 64'd4955519247014354852;
    12'd998: brom_out <= 64'd7738119443583029214;
    12'd2022: brom_out <= 64'd9080331558622478031;
    12'd22: brom_out <= 64'd4615809621887469834;
    12'd1046: brom_out <= 64'd7034035874218285317;
    12'd534: brom_out <= 64'd2050825072035144119;
    12'd1558: brom_out <= 64'd6150226684764233060;
    12'd278: brom_out <= 64'd39215274894679338;
    12'd1302: brom_out <= 64'd1392775048899804333;
    12'd790: brom_out <= 64'd1962272768984737496;
    12'd1814: brom_out <= 64'd6840536134827980412;
    12'd150: brom_out <= 64'd2316424835105438440;
    12'd1174: brom_out <= 64'd7255464637348812401;
    12'd662: brom_out <= 64'd5753795322756871121;
    12'd1686: brom_out <= 64'd4739227534138343988;
    12'd406: brom_out <= 64'd4480674382896232731;
    12'd1430: brom_out <= 64'd7860109258233506994;
    12'd918: brom_out <= 64'd8654722175613653276;
    12'd1942: brom_out <= 64'd3698113229434577276;
    12'd86: brom_out <= 64'd5761833653038383863;
    12'd1110: brom_out <= 64'd7649644688285296954;
    12'd598: brom_out <= 64'd5163048757488424028;
    12'd1622: brom_out <= 64'd280550462029244017;
    12'd342: brom_out <= 64'd2396874228472114740;
    12'd1366: brom_out <= 64'd367328239394980290;
    12'd854: brom_out <= 64'd1870367553472843855;
    12'd1878: brom_out <= 64'd242511422338012170;
    12'd214: brom_out <= 64'd7690852195393542907;
    12'd1238: brom_out <= 64'd6297789772157022780;
    12'd726: brom_out <= 64'd8943325242614027388;
    12'd1750: brom_out <= 64'd5788915943396697145;
    12'd470: brom_out <= 64'd2823654673579641862;
    12'd1494: brom_out <= 64'd2285701062711654789;
    12'd982: brom_out <= 64'd4735046624471887624;
    12'd2006: brom_out <= 64'd6703962736207848429;
    12'd54: brom_out <= 64'd437667873991410071;
    12'd1078: brom_out <= 64'd8941021957669153874;
    12'd566: brom_out <= 64'd5056679577221080592;
    12'd1590: brom_out <= 64'd7943456621955309555;
    12'd310: brom_out <= 64'd1663765558123988192;
    12'd1334: brom_out <= 64'd2197450412220039852;
    12'd822: brom_out <= 64'd6328044788619028811;
    12'd1846: brom_out <= 64'd5242800173554016477;
    12'd182: brom_out <= 64'd2051991327091467226;
    12'd1206: brom_out <= 64'd3566392214666874642;
    12'd694: brom_out <= 64'd3078044420483959468;
    12'd1718: brom_out <= 64'd2915851546318381008;
    12'd438: brom_out <= 64'd4973616575883620457;
    12'd1462: brom_out <= 64'd4590437479511182099;
    12'd950: brom_out <= 64'd1575596492305374553;
    12'd1974: brom_out <= 64'd7278311581654799448;
    12'd118: brom_out <= 64'd4255046251430904880;
    12'd1142: brom_out <= 64'd6014714335815937437;
    12'd630: brom_out <= 64'd5641268326478727432;
    12'd1654: brom_out <= 64'd3976255665346535912;
    12'd374: brom_out <= 64'd1523227976559640384;
    12'd1398: brom_out <= 64'd145908649510867226;
    12'd886: brom_out <= 64'd8191643213590331395;
    12'd1910: brom_out <= 64'd6676656787705972117;
    12'd246: brom_out <= 64'd838226266180407182;
    12'd1270: brom_out <= 64'd4147300013779743368;
    12'd758: brom_out <= 64'd4361527083377994653;
    12'd1782: brom_out <= 64'd7919187914793469944;
    12'd502: brom_out <= 64'd7725328103335519587;
    12'd1526: brom_out <= 64'd3130953281913181359;
    12'd1014: brom_out <= 64'd6038569734291399937;
    12'd2038: brom_out <= 64'd8186145541590340332;
    12'd14: brom_out <= 64'd8377422649175986985;
    12'd1038: brom_out <= 64'd4396018798804865849;
    12'd526: brom_out <= 64'd5298339161763062872;
    12'd1550: brom_out <= 64'd3031370596743080155;
    12'd270: brom_out <= 64'd772839773100063334;
    12'd1294: brom_out <= 64'd7106576547443304391;
    12'd782: brom_out <= 64'd8368352387789485495;
    12'd1806: brom_out <= 64'd4178694369519490509;
    12'd142: brom_out <= 64'd4118250476934667225;
    12'd1166: brom_out <= 64'd5668960288155274030;
    12'd654: brom_out <= 64'd6622650471528074404;
    12'd1678: brom_out <= 64'd4817909393282629696;
    12'd398: brom_out <= 64'd453516021392539197;
    12'd1422: brom_out <= 64'd6723432813723442718;
    12'd910: brom_out <= 64'd8804027098446734892;
    12'd1934: brom_out <= 64'd1882757962612426582;
    12'd78: brom_out <= 64'd2899615875029647480;
    12'd1102: brom_out <= 64'd9210839687198288177;
    12'd590: brom_out <= 64'd6180877422321376554;
    12'd1614: brom_out <= 64'd2226652841504127992;
    12'd334: brom_out <= 64'd1145275037428642328;
    12'd1358: brom_out <= 64'd2267277840274849562;
    12'd846: brom_out <= 64'd1986248922307912866;
    12'd1870: brom_out <= 64'd6322304445694945606;
    12'd206: brom_out <= 64'd4666975105442129532;
    12'd1230: brom_out <= 64'd7976502117851829149;
    12'd718: brom_out <= 64'd4385443872041495003;
    12'd1742: brom_out <= 64'd2564870828908612241;
    12'd462: brom_out <= 64'd8832127852899182441;
    12'd1486: brom_out <= 64'd2213631137681652193;
    12'd974: brom_out <= 64'd3122399872688598645;
    12'd1998: brom_out <= 64'd7569228676802102869;
    12'd46: brom_out <= 64'd8569730100285744993;
    12'd1070: brom_out <= 64'd7903746091327185660;
    12'd558: brom_out <= 64'd8659084273261581125;
    12'd1582: brom_out <= 64'd7661636433545697779;
    12'd302: brom_out <= 64'd5679245161077993970;
    12'd1326: brom_out <= 64'd2449958576690899108;
    12'd814: brom_out <= 64'd1269195536004574022;
    12'd1838: brom_out <= 64'd1447841990018008700;
    12'd174: brom_out <= 64'd5332325827108188102;
    12'd1198: brom_out <= 64'd8411339022167897455;
    12'd686: brom_out <= 64'd4717105437754674351;
    12'd1710: brom_out <= 64'd1292060914126343164;
    12'd430: brom_out <= 64'd7633783851459185362;
    12'd1454: brom_out <= 64'd309973352423096666;
    12'd942: brom_out <= 64'd1770807427320998317;
    12'd1966: brom_out <= 64'd8452824607548535710;
    12'd110: brom_out <= 64'd4414872346084808432;
    12'd1134: brom_out <= 64'd7826911971916988528;
    12'd622: brom_out <= 64'd234758437587011249;
    12'd1646: brom_out <= 64'd1144787620077612517;
    12'd366: brom_out <= 64'd4868519858037319455;
    12'd1390: brom_out <= 64'd2323588586179697296;
    12'd878: brom_out <= 64'd5022095663321251929;
    12'd1902: brom_out <= 64'd3131032845833922476;
    12'd238: brom_out <= 64'd9131483397025986172;
    12'd1262: brom_out <= 64'd3631295184904577614;
    12'd750: brom_out <= 64'd5571900938877394985;
    12'd1774: brom_out <= 64'd8150576788697059777;
    12'd494: brom_out <= 64'd4686751576350869864;
    12'd1518: brom_out <= 64'd7423219827873080903;
    12'd1006: brom_out <= 64'd6214632903940924813;
    12'd2030: brom_out <= 64'd2367595077715273251;
    12'd30: brom_out <= 64'd6118574647859303507;
    12'd1054: brom_out <= 64'd3858760292944247421;
    12'd542: brom_out <= 64'd1839144785420288440;
    12'd1566: brom_out <= 64'd4907547292263365345;
    12'd286: brom_out <= 64'd2615350370399979987;
    12'd1310: brom_out <= 64'd7271930591443660967;
    12'd798: brom_out <= 64'd6691738179524093988;
    12'd1822: brom_out <= 64'd6975474022730819773;
    12'd158: brom_out <= 64'd1817840973702651488;
    12'd1182: brom_out <= 64'd3375222894672577016;
    12'd670: brom_out <= 64'd2947366737269368820;
    12'd1694: brom_out <= 64'd1948091435642752956;
    12'd414: brom_out <= 64'd5140028477110672024;
    12'd1438: brom_out <= 64'd7172788441516230811;
    12'd926: brom_out <= 64'd8856614942545011767;
    12'd1950: brom_out <= 64'd1327034689155656339;
    12'd94: brom_out <= 64'd8469914002463831677;
    12'd1118: brom_out <= 64'd2146758214097748109;
    12'd606: brom_out <= 64'd8588335613155464482;
    12'd1630: brom_out <= 64'd317578861858216246;
    12'd350: brom_out <= 64'd2141294836449679462;
    12'd1374: brom_out <= 64'd8418770681392400674;
    12'd862: brom_out <= 64'd3513720992265299851;
    12'd1886: brom_out <= 64'd8399617655987284291;
    12'd222: brom_out <= 64'd2432371469911686242;
    12'd1246: brom_out <= 64'd8604033891536029454;
    12'd734: brom_out <= 64'd7837424891880392074;
    12'd1758: brom_out <= 64'd4686405902060845476;
    12'd478: brom_out <= 64'd6967909102360836955;
    12'd1502: brom_out <= 64'd3857651597088277268;
    12'd990: brom_out <= 64'd1834004577601037434;
    12'd2014: brom_out <= 64'd8282194139636476135;
    12'd62: brom_out <= 64'd7678547671088424856;
    12'd1086: brom_out <= 64'd2720286184019025751;
    12'd574: brom_out <= 64'd9012952791921640045;
    12'd1598: brom_out <= 64'd2141119197798094365;
    12'd318: brom_out <= 64'd3022986537941982063;
    12'd1342: brom_out <= 64'd4018445820304089225;
    12'd830: brom_out <= 64'd3518554950637655974;
    12'd1854: brom_out <= 64'd4340062858161126795;
    12'd190: brom_out <= 64'd8290294949532754385;
    12'd1214: brom_out <= 64'd7377937203894012946;
    12'd702: brom_out <= 64'd329797765029654054;
    12'd1726: brom_out <= 64'd7014388834507698157;
    12'd446: brom_out <= 64'd6987291732723720400;
    12'd1470: brom_out <= 64'd1664574738286193880;
    12'd958: brom_out <= 64'd5208572528313800398;
    12'd1982: brom_out <= 64'd7911339401561392797;
    12'd126: brom_out <= 64'd5187209805228830799;
    12'd1150: brom_out <= 64'd2094950622026922337;
    12'd638: brom_out <= 64'd2028205246324844013;
    12'd1662: brom_out <= 64'd8339080127670012014;
    12'd382: brom_out <= 64'd4524030704784542908;
    12'd1406: brom_out <= 64'd5544732514213129286;
    12'd894: brom_out <= 64'd4261169592821314574;
    12'd1918: brom_out <= 64'd4979449469273754225;
    12'd254: brom_out <= 64'd1956128207780189635;
    12'd1278: brom_out <= 64'd4026729170418869818;
    12'd766: brom_out <= 64'd5876647702261231319;
    12'd1790: brom_out <= 64'd398304142279976468;
    12'd510: brom_out <= 64'd4630776278738159906;
    12'd1534: brom_out <= 64'd3185152952275971112;
    12'd1022: brom_out <= 64'd8257506376334025193;
    12'd2046: brom_out <= 64'd5698772498710898262;
    12'd1: brom_out <= 64'd3410699927997700992;
    12'd1025: brom_out <= 64'd5129215985359186517;
    12'd513: brom_out <= 64'd6054184119640323055;
    12'd1537: brom_out <= 64'd8036011169461246502;
    12'd257: brom_out <= 64'd7134634440556594085;
    12'd1281: brom_out <= 64'd3042202103199590713;
    12'd769: brom_out <= 64'd4281242190677458415;
    12'd1793: brom_out <= 64'd5213930877604378225;
    12'd129: brom_out <= 64'd744370452723351798;
    12'd1153: brom_out <= 64'd386092701622236123;
    12'd641: brom_out <= 64'd1536404463035500281;
    12'd1665: brom_out <= 64'd3634367512595425146;
    12'd385: brom_out <= 64'd6470321026658955762;
    12'd1409: brom_out <= 64'd7247527117994054101;
    12'd897: brom_out <= 64'd5966322267827257001;
    12'd1921: brom_out <= 64'd8143790397219762868;
    12'd65: brom_out <= 64'd2548606593438851845;
    12'd1089: brom_out <= 64'd3842896822460231136;
    12'd577: brom_out <= 64'd7560481719955582125;
    12'd1601: brom_out <= 64'd4077854330096076199;
    12'd321: brom_out <= 64'd2524729693769219972;
    12'd1345: brom_out <= 64'd8864049892050671558;
    12'd833: brom_out <= 64'd4817445009517402390;
    12'd1857: brom_out <= 64'd7447202594453975344;
    12'd193: brom_out <= 64'd5467481028975156710;
    12'd1217: brom_out <= 64'd5274738861866299769;
    12'd705: brom_out <= 64'd5622958833092790840;
    12'd1729: brom_out <= 64'd6534274900636055338;
    12'd449: brom_out <= 64'd772485472146373328;
    12'd1473: brom_out <= 64'd189794809580270049;
    12'd961: brom_out <= 64'd3547010662611239126;
    12'd1985: brom_out <= 64'd5032432111932543760;
    12'd33: brom_out <= 64'd2256281196872481285;
    12'd1057: brom_out <= 64'd244042904533989192;
    12'd545: brom_out <= 64'd7081127620871813907;
    12'd1569: brom_out <= 64'd5045183220055932261;
    12'd289: brom_out <= 64'd155275333900253180;
    12'd1313: brom_out <= 64'd5068961430502894913;
    12'd801: brom_out <= 64'd6609966424554171950;
    12'd1825: brom_out <= 64'd8987443061574778656;
    12'd161: brom_out <= 64'd378592061626323514;
    12'd1185: brom_out <= 64'd8795660516396472524;
    12'd673: brom_out <= 64'd4904003744551651835;
    12'd1697: brom_out <= 64'd6139101682900360503;
    12'd417: brom_out <= 64'd2682034885057011637;
    12'd1441: brom_out <= 64'd3477251427531362048;
    12'd929: brom_out <= 64'd7073132918750649160;
    12'd1953: brom_out <= 64'd2334160254732771581;
    12'd97: brom_out <= 64'd2888862071876983052;
    12'd1121: brom_out <= 64'd2156941117628995192;
    12'd609: brom_out <= 64'd5073469937111083807;
    12'd1633: brom_out <= 64'd4840479360880356651;
    12'd353: brom_out <= 64'd5421857412712885675;
    12'd1377: brom_out <= 64'd162811161267629503;
    12'd865: brom_out <= 64'd5646027969675254732;
    12'd1889: brom_out <= 64'd755640484730109350;
    12'd225: brom_out <= 64'd2826479692684020797;
    12'd1249: brom_out <= 64'd219379608293825313;
    12'd737: brom_out <= 64'd764974623599952144;
    12'd1761: brom_out <= 64'd214719891515706016;
    12'd481: brom_out <= 64'd6589512973569282125;
    12'd1505: brom_out <= 64'd1934857541461099950;
    12'd993: brom_out <= 64'd7177314716649923316;
    12'd2017: brom_out <= 64'd7922313050019057439;
    12'd17: brom_out <= 64'd3362845476240585630;
    12'd1041: brom_out <= 64'd4404677075369256989;
    12'd529: brom_out <= 64'd2418333291631172466;
    12'd1553: brom_out <= 64'd6230802514162268134;
    12'd273: brom_out <= 64'd3341668352136705219;
    12'd1297: brom_out <= 64'd8956370168834558428;
    12'd785: brom_out <= 64'd7608656401006491194;
    12'd1809: brom_out <= 64'd698708485609276696;
    12'd145: brom_out <= 64'd3058030583995206520;
    12'd1169: brom_out <= 64'd353110664605704442;
    12'd657: brom_out <= 64'd3017120554102128340;
    12'd1681: brom_out <= 64'd5103733993327281237;
    12'd401: brom_out <= 64'd2741677917677613231;
    12'd1425: brom_out <= 64'd8662664786796030150;
    12'd913: brom_out <= 64'd763839710936525575;
    12'd1937: brom_out <= 64'd347979942635009334;
    12'd81: brom_out <= 64'd7976504752654974117;
    12'd1105: brom_out <= 64'd3436462466961844858;
    12'd593: brom_out <= 64'd4429449008218948808;
    12'd1617: brom_out <= 64'd2658082230673248031;
    12'd337: brom_out <= 64'd7185619194359065362;
    12'd1361: brom_out <= 64'd1114116847695536049;
    12'd849: brom_out <= 64'd884137179653819607;
    12'd1873: brom_out <= 64'd5065067130629118737;
    12'd209: brom_out <= 64'd8393585351321635411;
    12'd1233: brom_out <= 64'd7090807160606196052;
    12'd721: brom_out <= 64'd6410485094202897752;
    12'd1745: brom_out <= 64'd9022101888677434117;
    12'd465: brom_out <= 64'd1589614425957732699;
    12'd1489: brom_out <= 64'd6013752395227127263;
    12'd977: brom_out <= 64'd3386135057788622513;
    12'd2001: brom_out <= 64'd1330478846821969397;
    12'd49: brom_out <= 64'd386281610427438192;
    12'd1073: brom_out <= 64'd2035588011496638896;
    12'd561: brom_out <= 64'd4232540739601334965;
    12'd1585: brom_out <= 64'd1859092738452818058;
    12'd305: brom_out <= 64'd6645577682609730772;
    12'd1329: brom_out <= 64'd983596768654482029;
    12'd817: brom_out <= 64'd2156960173702089180;
    12'd1841: brom_out <= 64'd1429662614925885796;
    12'd177: brom_out <= 64'd2864911663037216672;
    12'd1201: brom_out <= 64'd5334612837580195271;
    12'd689: brom_out <= 64'd4228541773534977716;
    12'd1713: brom_out <= 64'd3892775677548530090;
    12'd433: brom_out <= 64'd5044810319583755777;
    12'd1457: brom_out <= 64'd7352579042178488139;
    12'd945: brom_out <= 64'd1952516211385548365;
    12'd1969: brom_out <= 64'd5262043117036187744;
    12'd113: brom_out <= 64'd4738275030069272353;
    12'd1137: brom_out <= 64'd8415750935695247922;
    12'd625: brom_out <= 64'd4325481024329050713;
    12'd1649: brom_out <= 64'd7746766013427248385;
    12'd369: brom_out <= 64'd2556972555839883886;
    12'd1393: brom_out <= 64'd6044588417436356179;
    12'd881: brom_out <= 64'd3666634855840044384;
    12'd1905: brom_out <= 64'd1611916591103368969;
    12'd241: brom_out <= 64'd4992072784223513734;
    12'd1265: brom_out <= 64'd3829684802947366251;
    12'd753: brom_out <= 64'd6613926690929773980;
    12'd1777: brom_out <= 64'd5622262333701922490;
    12'd497: brom_out <= 64'd2811982284434465810;
    12'd1521: brom_out <= 64'd4967992377336504914;
    12'd1009: brom_out <= 64'd997335904832336470;
    12'd2033: brom_out <= 64'd4820986686989856162;
    12'd9: brom_out <= 64'd765633873015113116;
    12'd1033: brom_out <= 64'd7788210691976825999;
    12'd521: brom_out <= 64'd6235145204509423075;
    12'd1545: brom_out <= 64'd1118292230605154455;
    12'd265: brom_out <= 64'd6297397295888024961;
    12'd1289: brom_out <= 64'd5917236050195909530;
    12'd777: brom_out <= 64'd7377440782932470849;
    12'd1801: brom_out <= 64'd139707927547171638;
    12'd137: brom_out <= 64'd4144450591698584079;
    12'd1161: brom_out <= 64'd9070945006014315493;
    12'd649: brom_out <= 64'd4795769251779777619;
    12'd1673: brom_out <= 64'd3342253550284462446;
    12'd393: brom_out <= 64'd5441354093845414231;
    12'd1417: brom_out <= 64'd6918683828302718739;
    12'd905: brom_out <= 64'd734568655330607842;
    12'd1929: brom_out <= 64'd7857302122066421647;
    12'd73: brom_out <= 64'd3145931349312735151;
    12'd1097: brom_out <= 64'd8424370584387910975;
    12'd585: brom_out <= 64'd222811142323919754;
    12'd1609: brom_out <= 64'd7574831232213709396;
    12'd329: brom_out <= 64'd8043393289914459292;
    12'd1353: brom_out <= 64'd7244116446129534888;
    12'd841: brom_out <= 64'd5017580708797525693;
    12'd1865: brom_out <= 64'd6706908070502136570;
    12'd201: brom_out <= 64'd6711532558695792766;
    12'd1225: brom_out <= 64'd8975566828816296230;
    12'd713: brom_out <= 64'd9186619957940342983;
    12'd1737: brom_out <= 64'd6575585304828318751;
    12'd457: brom_out <= 64'd8454482646563058332;
    12'd1481: brom_out <= 64'd6033474465198015463;
    12'd969: brom_out <= 64'd7175151278796593227;
    12'd1993: brom_out <= 64'd2486042518374802962;
    12'd41: brom_out <= 64'd6198065040356620108;
    12'd1065: brom_out <= 64'd8612567367455566604;
    12'd553: brom_out <= 64'd8848185420485894564;
    12'd1577: brom_out <= 64'd4191997763519057770;
    12'd297: brom_out <= 64'd2139183688024244662;
    12'd1321: brom_out <= 64'd2416292409822388515;
    12'd809: brom_out <= 64'd262231450558211361;
    12'd1833: brom_out <= 64'd4587030516195245229;
    12'd169: brom_out <= 64'd1415022612836804245;
    12'd1193: brom_out <= 64'd3995462545347869825;
    12'd681: brom_out <= 64'd7666496919135739619;
    12'd1705: brom_out <= 64'd3616245215788926208;
    12'd425: brom_out <= 64'd3402060265689055646;
    12'd1449: brom_out <= 64'd8241718962591948447;
    12'd937: brom_out <= 64'd4573518681633497875;
    12'd1961: brom_out <= 64'd588418346038461962;
    12'd105: brom_out <= 64'd4387570214710289221;
    12'd1129: brom_out <= 64'd5478727957299769295;
    12'd617: brom_out <= 64'd8357119822637878344;
    12'd1641: brom_out <= 64'd603953902387193508;
    12'd361: brom_out <= 64'd6543748061310240720;
    12'd1385: brom_out <= 64'd7668686831057436985;
    12'd873: brom_out <= 64'd3935686344822117526;
    12'd1897: brom_out <= 64'd6181451780242161625;
    12'd233: brom_out <= 64'd409924620725067559;
    12'd1257: brom_out <= 64'd7892948909074176925;
    12'd745: brom_out <= 64'd6226526169594591809;
    12'd1769: brom_out <= 64'd9134180865229835759;
    12'd489: brom_out <= 64'd4490148815910336990;
    12'd1513: brom_out <= 64'd2355439580988530149;
    12'd1001: brom_out <= 64'd6518635118472409845;
    12'd2025: brom_out <= 64'd51936672487212441;
    12'd25: brom_out <= 64'd6715985458946590128;
    12'd1049: brom_out <= 64'd5762672832480805366;
    12'd537: brom_out <= 64'd2995687659634637462;
    12'd1561: brom_out <= 64'd7461219876635110075;
    12'd281: brom_out <= 64'd7183447847060170764;
    12'd1305: brom_out <= 64'd1183708660053992021;
    12'd793: brom_out <= 64'd5777835500516375970;
    12'd1817: brom_out <= 64'd5095646658923524735;
    12'd153: brom_out <= 64'd3113727683625837877;
    12'd1177: brom_out <= 64'd2523123097999550009;
    12'd665: brom_out <= 64'd7142186205919208875;
    12'd1689: brom_out <= 64'd9217750718102413769;
    12'd409: brom_out <= 64'd1657391714823220364;
    12'd1433: brom_out <= 64'd3134034012266112081;
    12'd921: brom_out <= 64'd8791253981502320058;
    12'd1945: brom_out <= 64'd4661856834147524101;
    12'd89: brom_out <= 64'd4869054365853473205;
    12'd1113: brom_out <= 64'd282601018708895118;
    12'd601: brom_out <= 64'd6393795207000798995;
    12'd1625: brom_out <= 64'd7025885032724338522;
    12'd345: brom_out <= 64'd4568626412972067498;
    12'd1369: brom_out <= 64'd2863468293897413688;
    12'd857: brom_out <= 64'd4813342945543862763;
    12'd1881: brom_out <= 64'd2716283261879775205;
    12'd217: brom_out <= 64'd3010181431159388657;
    12'd1241: brom_out <= 64'd955620117667129746;
    12'd729: brom_out <= 64'd133811528865334890;
    12'd1753: brom_out <= 64'd1833025850275574712;
    12'd473: brom_out <= 64'd7876920601219670377;
    12'd1497: brom_out <= 64'd6527564409825216632;
    12'd985: brom_out <= 64'd1514716156703592623;
    12'd2009: brom_out <= 64'd4985122398795428546;
    12'd57: brom_out <= 64'd6345337778311606873;
    12'd1081: brom_out <= 64'd3401727224945347906;
    12'd569: brom_out <= 64'd47457376937832185;
    12'd1593: brom_out <= 64'd852557670474817786;
    12'd313: brom_out <= 64'd8123831902889627067;
    12'd1337: brom_out <= 64'd2384224833012558450;
    12'd825: brom_out <= 64'd2796841718743354108;
    12'd1849: brom_out <= 64'd8015393524551084254;
    12'd185: brom_out <= 64'd5237617555609021497;
    12'd1209: brom_out <= 64'd5012862545847756521;
    12'd697: brom_out <= 64'd6366523862546675874;
    12'd1721: brom_out <= 64'd3778417854489625020;
    12'd441: brom_out <= 64'd7188215029319270896;
    12'd1465: brom_out <= 64'd6695490825212130486;
    12'd953: brom_out <= 64'd8903646571445642590;
    12'd1977: brom_out <= 64'd3058024851622871963;
    12'd121: brom_out <= 64'd2537688559670774442;
    12'd1145: brom_out <= 64'd886809128212118598;
    12'd633: brom_out <= 64'd7697594985778228047;
    12'd1657: brom_out <= 64'd4395955890441811094;
    12'd377: brom_out <= 64'd100480137207823859;
    12'd1401: brom_out <= 64'd110551151910388577;
    12'd889: brom_out <= 64'd3189663103820318230;
    12'd1913: brom_out <= 64'd2379296037912008850;
    12'd249: brom_out <= 64'd2763047856760583059;
    12'd1273: brom_out <= 64'd6756397676980789867;
    12'd761: brom_out <= 64'd7207388653722405316;
    12'd1785: brom_out <= 64'd1943133841497291102;
    12'd505: brom_out <= 64'd2552637224532115932;
    12'd1529: brom_out <= 64'd6598765433084769229;
    12'd1017: brom_out <= 64'd2320923143671569896;
    12'd2041: brom_out <= 64'd5556671996955451950;
    12'd5: brom_out <= 64'd6763758159452639774;
    12'd1029: brom_out <= 64'd2267375919945251521;
    12'd517: brom_out <= 64'd454590519805025044;
    12'd1541: brom_out <= 64'd6304263996515549886;
    12'd261: brom_out <= 64'd9197007911222417389;
    12'd1285: brom_out <= 64'd2377243651087003666;
    12'd773: brom_out <= 64'd6143431748742725020;
    12'd1797: brom_out <= 64'd5354215831080117776;
    12'd133: brom_out <= 64'd6016428244618191862;
    12'd1157: brom_out <= 64'd4382417857856181174;
    12'd645: brom_out <= 64'd7751899648531048175;
    12'd1669: brom_out <= 64'd2630294209519613088;
    12'd389: brom_out <= 64'd1501378395168039326;
    12'd1413: brom_out <= 64'd8551983914694877356;
    12'd901: brom_out <= 64'd2906457744329251012;
    12'd1925: brom_out <= 64'd5286915306002180265;
    12'd69: brom_out <= 64'd1947002332183469414;
    12'd1093: brom_out <= 64'd96863724318406758;
    12'd581: brom_out <= 64'd2897620933911650343;
    12'd1605: brom_out <= 64'd4955839328155437349;
    12'd325: brom_out <= 64'd7481124282822080413;
    12'd1349: brom_out <= 64'd7020449510915630462;
    12'd837: brom_out <= 64'd508780516872826234;
    12'd1861: brom_out <= 64'd8016279939582392242;
    12'd197: brom_out <= 64'd2595662895600887742;
    12'd1221: brom_out <= 64'd6466645302876820970;
    12'd709: brom_out <= 64'd5711044082124335681;
    12'd1733: brom_out <= 64'd1232589470396273160;
    12'd453: brom_out <= 64'd2672804684031921286;
    12'd1477: brom_out <= 64'd2366301485405412450;
    12'd965: brom_out <= 64'd2110442893422689640;
    12'd1989: brom_out <= 64'd1718577144632118127;
    12'd37: brom_out <= 64'd4813944553649371399;
    12'd1061: brom_out <= 64'd4255745979415696947;
    12'd549: brom_out <= 64'd4023116666530304294;
    12'd1573: brom_out <= 64'd3357048858130187252;
    12'd293: brom_out <= 64'd1600525449816895321;
    12'd1317: brom_out <= 64'd1300018304757311460;
    12'd805: brom_out <= 64'd2181414353711885500;
    12'd1829: brom_out <= 64'd3950462616828770811;
    12'd165: brom_out <= 64'd1946463679777770624;
    12'd1189: brom_out <= 64'd4547618201573256410;
    12'd677: brom_out <= 64'd7238012484886626569;
    12'd1701: brom_out <= 64'd536380155698109790;
    12'd421: brom_out <= 64'd8270909668692229778;
    12'd1445: brom_out <= 64'd3811108364812692601;
    12'd933: brom_out <= 64'd6648757142176170015;
    12'd1957: brom_out <= 64'd5629290568836098156;
    12'd101: brom_out <= 64'd2178058660755934531;
    12'd1125: brom_out <= 64'd1126887764375740643;
    12'd613: brom_out <= 64'd1742705753673391143;
    12'd1637: brom_out <= 64'd6765134044717755623;
    12'd357: brom_out <= 64'd9212280164341746403;
    12'd1381: brom_out <= 64'd1433093515373313065;
    12'd869: brom_out <= 64'd7877777968461631808;
    12'd1893: brom_out <= 64'd8785867091986638617;
    12'd229: brom_out <= 64'd485061594959071822;
    12'd1253: brom_out <= 64'd989361657948442110;
    12'd741: brom_out <= 64'd2076728825140822847;
    12'd1765: brom_out <= 64'd3456130262014008515;
    12'd485: brom_out <= 64'd8278479492455693015;
    12'd1509: brom_out <= 64'd9195646169382126030;
    12'd997: brom_out <= 64'd5212168841016919149;
    12'd2021: brom_out <= 64'd9128090719146323475;
    12'd21: brom_out <= 64'd8164891973823639038;
    12'd1045: brom_out <= 64'd3746430640008993009;
    12'd533: brom_out <= 64'd5370605519979511464;
    12'd1557: brom_out <= 64'd7627180408796406893;
    12'd277: brom_out <= 64'd5555140140749937950;
    12'd1301: brom_out <= 64'd7404484841390992291;
    12'd789: brom_out <= 64'd7454066665886887296;
    12'd1813: brom_out <= 64'd1162336423194039634;
    12'd149: brom_out <= 64'd6781156493805473184;
    12'd1173: brom_out <= 64'd4194093989176669544;
    12'd661: brom_out <= 64'd4838827599606243518;
    12'd1685: brom_out <= 64'd2155237171088034080;
    12'd405: brom_out <= 64'd1238087211225650716;
    12'd1429: brom_out <= 64'd2685797616310619352;
    12'd917: brom_out <= 64'd1843312381298496268;
    12'd1941: brom_out <= 64'd2162964054538971540;
    12'd85: brom_out <= 64'd1894954218249665392;
    12'd1109: brom_out <= 64'd6484383960926813681;
    12'd597: brom_out <= 64'd7646724549737265499;
    12'd1621: brom_out <= 64'd6205849589163236816;
    12'd341: brom_out <= 64'd1301636535530801539;
    12'd1365: brom_out <= 64'd5282390222647191044;
    12'd853: brom_out <= 64'd2771334574021323382;
    12'd1877: brom_out <= 64'd2385017937900592304;
    12'd213: brom_out <= 64'd1151378716197177552;
    12'd1237: brom_out <= 64'd709914170400347798;
    12'd725: brom_out <= 64'd5274592101237787712;
    12'd1749: brom_out <= 64'd8291454664421844925;
    12'd469: brom_out <= 64'd7662747679479933417;
    12'd1493: brom_out <= 64'd7481296381304816625;
    12'd981: brom_out <= 64'd414905064980978750;
    12'd2005: brom_out <= 64'd6111286953235601862;
    12'd53: brom_out <= 64'd7624179653698414196;
    12'd1077: brom_out <= 64'd3154230262077045121;
    12'd565: brom_out <= 64'd3988697203834155060;
    12'd1589: brom_out <= 64'd8542379982640788350;
    12'd309: brom_out <= 64'd6544569414691682489;
    12'd1333: brom_out <= 64'd2183199595637029406;
    12'd821: brom_out <= 64'd4670201655156419723;
    12'd1845: brom_out <= 64'd5498459411109788068;
    12'd181: brom_out <= 64'd4278858494259842183;
    12'd1205: brom_out <= 64'd7796442270140558508;
    12'd693: brom_out <= 64'd4857978139238569870;
    12'd1717: brom_out <= 64'd6399210596466476392;
    12'd437: brom_out <= 64'd6096366000398327739;
    12'd1461: brom_out <= 64'd1867571504953480770;
    12'd949: brom_out <= 64'd3412217070080433702;
    12'd1973: brom_out <= 64'd4577353689341769269;
    12'd117: brom_out <= 64'd3008075931742456305;
    12'd1141: brom_out <= 64'd876318092677120142;
    12'd629: brom_out <= 64'd1717951383164415823;
    12'd1653: brom_out <= 64'd3169734437867057239;
    12'd373: brom_out <= 64'd4767362740579418704;
    12'd1397: brom_out <= 64'd5650772903320476912;
    12'd885: brom_out <= 64'd5653087238811240759;
    12'd1909: brom_out <= 64'd1189621726592624294;
    12'd245: brom_out <= 64'd9221845814575141125;
    12'd1269: brom_out <= 64'd4660090867314689002;
    12'd757: brom_out <= 64'd2242075921938682459;
    12'd1781: brom_out <= 64'd3116024623734582454;
    12'd501: brom_out <= 64'd3036549354902120193;
    12'd1525: brom_out <= 64'd5042277015269219313;
    12'd1013: brom_out <= 64'd3484131572223489484;
    12'd2037: brom_out <= 64'd961913442728646227;
    12'd13: brom_out <= 64'd1308543301457948090;
    12'd1037: brom_out <= 64'd3637382950058536861;
    12'd525: brom_out <= 64'd1393749877433722763;
    12'd1549: brom_out <= 64'd537819627866893722;
    12'd269: brom_out <= 64'd6447255846682879893;
    12'd1293: brom_out <= 64'd8786731256157126405;
    12'd781: brom_out <= 64'd3997949459943286754;
    12'd1805: brom_out <= 64'd8324077327553852513;
    12'd141: brom_out <= 64'd7394755339662913294;
    12'd1165: brom_out <= 64'd4673703781571774967;
    12'd653: brom_out <= 64'd1728666539874811802;
    12'd1677: brom_out <= 64'd4057021711048425673;
    12'd397: brom_out <= 64'd566944775070236995;
    12'd1421: brom_out <= 64'd2547651610572949376;
    12'd909: brom_out <= 64'd2329726160784570819;
    12'd1933: brom_out <= 64'd1161862294465578057;
    12'd77: brom_out <= 64'd4644587485367466700;
    12'd1101: brom_out <= 64'd5294971316032015895;
    12'd589: brom_out <= 64'd5912831972142402456;
    12'd1613: brom_out <= 64'd5795447197771939000;
    12'd333: brom_out <= 64'd1686606374247730404;
    12'd1357: brom_out <= 64'd6092744959824246525;
    12'd845: brom_out <= 64'd1618740323245231299;
    12'd1869: brom_out <= 64'd8598342625683728299;
    12'd205: brom_out <= 64'd8817740569999643205;
    12'd1229: brom_out <= 64'd6960470765855428832;
    12'd717: brom_out <= 64'd2337429885856105847;
    12'd1741: brom_out <= 64'd5179217325409368865;
    12'd461: brom_out <= 64'd6106183392065786101;
    12'd1485: brom_out <= 64'd4024635328045370383;
    12'd973: brom_out <= 64'd6235292595162042788;
    12'd1997: brom_out <= 64'd6868627029504454320;
    12'd45: brom_out <= 64'd3756196661099655504;
    12'd1069: brom_out <= 64'd8553381754481976676;
    12'd557: brom_out <= 64'd4862932399326851702;
    12'd1581: brom_out <= 64'd2657217402772260763;
    12'd301: brom_out <= 64'd4523637763894961641;
    12'd1325: brom_out <= 64'd3292349049063742778;
    12'd813: brom_out <= 64'd9155970337107209825;
    12'd1837: brom_out <= 64'd3997725441927781364;
    12'd173: brom_out <= 64'd4740834202485229233;
    12'd1197: brom_out <= 64'd4066382155101871051;
    12'd685: brom_out <= 64'd508271619034446786;
    12'd1709: brom_out <= 64'd7401485280983992861;
    12'd429: brom_out <= 64'd5082132714401984683;
    12'd1453: brom_out <= 64'd333880186367592003;
    12'd941: brom_out <= 64'd5446865046789948513;
    12'd1965: brom_out <= 64'd2725414062112306281;
    12'd109: brom_out <= 64'd1248372373386200542;
    12'd1133: brom_out <= 64'd1119335065523703938;
    12'd621: brom_out <= 64'd7840124210205868861;
    12'd1645: brom_out <= 64'd3023524884400278775;
    12'd365: brom_out <= 64'd2736243621131921998;
    12'd1389: brom_out <= 64'd3539469165500234284;
    12'd877: brom_out <= 64'd1888290614954743033;
    12'd1901: brom_out <= 64'd7520330660356266028;
    12'd237: brom_out <= 64'd6863887312817181582;
    12'd1261: brom_out <= 64'd6398295448536016830;
    12'd749: brom_out <= 64'd1592524290669994207;
    12'd1773: brom_out <= 64'd5910759767512541250;
    12'd493: brom_out <= 64'd3830971498294533116;
    12'd1517: brom_out <= 64'd8956726076603480703;
    12'd1005: brom_out <= 64'd2589999426439265259;
    12'd2029: brom_out <= 64'd4970849700277405618;
    12'd29: brom_out <= 64'd5273329109373150975;
    12'd1053: brom_out <= 64'd7460628603806863746;
    12'd541: brom_out <= 64'd434031393225567768;
    12'd1565: brom_out <= 64'd8465546254545831686;
    12'd285: brom_out <= 64'd9078993651166531175;
    12'd1309: brom_out <= 64'd7807690460766985086;
    12'd797: brom_out <= 64'd8652975144754354580;
    12'd1821: brom_out <= 64'd1085102489027133340;
    12'd157: brom_out <= 64'd2743669863121200377;
    12'd1181: brom_out <= 64'd4467581496101227334;
    12'd669: brom_out <= 64'd3876556978203189868;
    12'd1693: brom_out <= 64'd4685721143967180157;
    12'd413: brom_out <= 64'd385686628599757307;
    12'd1437: brom_out <= 64'd2598484606631636222;
    12'd925: brom_out <= 64'd3535939462128378156;
    12'd1949: brom_out <= 64'd2577772307257209845;
    12'd93: brom_out <= 64'd946158067222968651;
    12'd1117: brom_out <= 64'd928066452629839385;
    12'd605: brom_out <= 64'd5206734552224755013;
    12'd1629: brom_out <= 64'd4014372500035666136;
    12'd349: brom_out <= 64'd2891611787780236417;
    12'd1373: brom_out <= 64'd2585495344379534056;
    12'd861: brom_out <= 64'd3338220124400918038;
    12'd1885: brom_out <= 64'd2576743551182428740;
    12'd221: brom_out <= 64'd8323498142012160010;
    12'd1245: brom_out <= 64'd4804504980610246604;
    12'd733: brom_out <= 64'd5684247906257495894;
    12'd1757: brom_out <= 64'd7951156483706292038;
    12'd477: brom_out <= 64'd2820663287170928640;
    12'd1501: brom_out <= 64'd5098869993716106906;
    12'd989: brom_out <= 64'd8866095157257406445;
    12'd2013: brom_out <= 64'd2660027230730544837;
    12'd61: brom_out <= 64'd1347697413910003923;
    12'd1085: brom_out <= 64'd2712792922253887919;
    12'd573: brom_out <= 64'd4376874011134652106;
    12'd1597: brom_out <= 64'd5396208835915368384;
    12'd317: brom_out <= 64'd7105200227530783706;
    12'd1341: brom_out <= 64'd3728375885890433547;
    12'd829: brom_out <= 64'd132470796801485904;
    12'd1853: brom_out <= 64'd3570793125845813024;
    12'd189: brom_out <= 64'd4908524226076483463;
    12'd1213: brom_out <= 64'd6302668669512474796;
    12'd701: brom_out <= 64'd1714417639468662926;
    12'd1725: brom_out <= 64'd1519611810510721602;
    12'd445: brom_out <= 64'd8839802895180069702;
    12'd1469: brom_out <= 64'd3044785443284390797;
    12'd957: brom_out <= 64'd3664031833482737832;
    12'd1981: brom_out <= 64'd8963319392399776246;
    12'd125: brom_out <= 64'd4480805174170202207;
    12'd1149: brom_out <= 64'd333389965294045693;
    12'd637: brom_out <= 64'd3741893797201556249;
    12'd1661: brom_out <= 64'd2000208331708224068;
    12'd381: brom_out <= 64'd7942507821398558532;
    12'd1405: brom_out <= 64'd6637586715306416768;
    12'd893: brom_out <= 64'd3321211816430529043;
    12'd1917: brom_out <= 64'd6308962713817541263;
    12'd253: brom_out <= 64'd6388259551719657978;
    12'd1277: brom_out <= 64'd1562593397733019041;
    12'd765: brom_out <= 64'd6219067382595841970;
    12'd1789: brom_out <= 64'd4841428800401574405;
    12'd509: brom_out <= 64'd3450684051664931847;
    12'd1533: brom_out <= 64'd574337591279463189;
    12'd1021: brom_out <= 64'd4361850440264709726;
    12'd2045: brom_out <= 64'd1440985375463933246;
    12'd3: brom_out <= 64'd3861962373613601910;
    12'd1027: brom_out <= 64'd4162209495553610418;
    12'd515: brom_out <= 64'd8043781972276579395;
    12'd1539: brom_out <= 64'd1340559018494124164;
    12'd259: brom_out <= 64'd3107882050279402743;
    12'd1283: brom_out <= 64'd7159694058507751872;
    12'd771: brom_out <= 64'd4005162996496124928;
    12'd1795: brom_out <= 64'd8529786556497506513;
    12'd131: brom_out <= 64'd1878779880994978994;
    12'd1155: brom_out <= 64'd5998107129159023210;
    12'd643: brom_out <= 64'd6012561626455134523;
    12'd1667: brom_out <= 64'd7471063379806895040;
    12'd387: brom_out <= 64'd2048632887949724958;
    12'd1411: brom_out <= 64'd3289993698217648619;
    12'd899: brom_out <= 64'd6442436536170659884;
    12'd1923: brom_out <= 64'd7317451652887540786;
    12'd67: brom_out <= 64'd1514048392223859021;
    12'd1091: brom_out <= 64'd1203672178180575298;
    12'd579: brom_out <= 64'd6380902013505704791;
    12'd1603: brom_out <= 64'd7430662062095694115;
    12'd323: brom_out <= 64'd5782810937935678862;
    12'd1347: brom_out <= 64'd2262139037550279899;
    12'd835: brom_out <= 64'd8305495959405484792;
    12'd1859: brom_out <= 64'd6490070968946649227;
    12'd195: brom_out <= 64'd2401026282272167012;
    12'd1219: brom_out <= 64'd5545997593461576288;
    12'd707: brom_out <= 64'd2666954462262670696;
    12'd1731: brom_out <= 64'd987669974730382046;
    12'd451: brom_out <= 64'd6458515334846772263;
    12'd1475: brom_out <= 64'd7249378466214688806;
    12'd963: brom_out <= 64'd5516671091365828465;
    12'd1987: brom_out <= 64'd8999967320369276511;
    12'd35: brom_out <= 64'd6062736565148073825;
    12'd1059: brom_out <= 64'd1608365741208693577;
    12'd547: brom_out <= 64'd7654152496553449131;
    12'd1571: brom_out <= 64'd4133493835850339168;
    12'd291: brom_out <= 64'd1585748934512571741;
    12'd1315: brom_out <= 64'd6612420970902801975;
    12'd803: brom_out <= 64'd454280960792274896;
    12'd1827: brom_out <= 64'd8497367263149911233;
    12'd163: brom_out <= 64'd5353640366896974923;
    12'd1187: brom_out <= 64'd6206358084041665071;
    12'd675: brom_out <= 64'd5272219219689335945;
    12'd1699: brom_out <= 64'd3803110647467949217;
    12'd419: brom_out <= 64'd1295390929475635113;
    12'd1443: brom_out <= 64'd4153998133878397451;
    12'd931: brom_out <= 64'd6620879955184290310;
    12'd1955: brom_out <= 64'd8754621773751208831;
    12'd99: brom_out <= 64'd2657155576256827462;
    12'd1123: brom_out <= 64'd8834017661859685034;
    12'd611: brom_out <= 64'd6843337341430130824;
    12'd1635: brom_out <= 64'd763353675495114124;
    12'd355: brom_out <= 64'd1133977356953084162;
    12'd1379: brom_out <= 64'd236770855711589184;
    12'd867: brom_out <= 64'd133065795425889836;
    12'd1891: brom_out <= 64'd2547546770525996332;
    12'd227: brom_out <= 64'd8686764207920541366;
    12'd1251: brom_out <= 64'd8237006339815446938;
    12'd739: brom_out <= 64'd8525414979588871296;
    12'd1763: brom_out <= 64'd2028388940891580996;
    12'd483: brom_out <= 64'd6576516027170948233;
    12'd1507: brom_out <= 64'd7339842136519118186;
    12'd995: brom_out <= 64'd6788808489126092282;
    12'd2019: brom_out <= 64'd9040689692862409764;
    12'd19: brom_out <= 64'd6708106808539775657;
    12'd1043: brom_out <= 64'd5205848358505084751;
    12'd531: brom_out <= 64'd3878767790153268931;
    12'd1555: brom_out <= 64'd796613256859496714;
    12'd275: brom_out <= 64'd7472637614049421408;
    12'd1299: brom_out <= 64'd1889553700543734703;
    12'd787: brom_out <= 64'd5854390915714537768;
    12'd1811: brom_out <= 64'd5788872167869932214;
    12'd147: brom_out <= 64'd907092075277997974;
    12'd1171: brom_out <= 64'd1839345025779015562;
    12'd659: brom_out <= 64'd6443072913543794285;
    12'd1683: brom_out <= 64'd5275675377974681218;
    12'd403: brom_out <= 64'd428290208011211366;
    12'd1427: brom_out <= 64'd5569321792001207118;
    12'd915: brom_out <= 64'd1977776347539890920;
    12'd1939: brom_out <= 64'd3135574699227801344;
    12'd83: brom_out <= 64'd689809073466025184;
    12'd1107: brom_out <= 64'd5624842936299281778;
    12'd595: brom_out <= 64'd5307440016266556877;
    12'd1619: brom_out <= 64'd8493599686472256014;
    12'd339: brom_out <= 64'd2227351510237238216;
    12'd1363: brom_out <= 64'd6377822362516206160;
    12'd851: brom_out <= 64'd898522998319472068;
    12'd1875: brom_out <= 64'd489770987855749055;
    12'd211: brom_out <= 64'd4043139279432890725;
    12'd1235: brom_out <= 64'd1876332191965133731;
    12'd723: brom_out <= 64'd5506819904638189904;
    12'd1747: brom_out <= 64'd5886621447526459673;
    12'd467: brom_out <= 64'd2808072814625355654;
    12'd1491: brom_out <= 64'd6516876726075941552;
    12'd979: brom_out <= 64'd1088097907932407751;
    12'd2003: brom_out <= 64'd5656721139433476677;
    12'd51: brom_out <= 64'd8944778841024587087;
    12'd1075: brom_out <= 64'd4893012051863450219;
    12'd563: brom_out <= 64'd4221070846363861203;
    12'd1587: brom_out <= 64'd3655024687870693466;
    12'd307: brom_out <= 64'd1652845580397658846;
    12'd1331: brom_out <= 64'd3994442180932799364;
    12'd819: brom_out <= 64'd4340151557824599919;
    12'd1843: brom_out <= 64'd6911465924675166044;
    12'd179: brom_out <= 64'd2914506150870709118;
    12'd1203: brom_out <= 64'd2222396136948961372;
    12'd691: brom_out <= 64'd6398233032526050184;
    12'd1715: brom_out <= 64'd8254701148114518467;
    12'd435: brom_out <= 64'd8629791111789113940;
    12'd1459: brom_out <= 64'd8971031896351058404;
    12'd947: brom_out <= 64'd1119603175546581820;
    12'd1971: brom_out <= 64'd5082461315959087042;
    12'd115: brom_out <= 64'd835265111212787639;
    12'd1139: brom_out <= 64'd8864546665859549780;
    12'd627: brom_out <= 64'd6349714072416716427;
    12'd1651: brom_out <= 64'd6191860356230181438;
    12'd371: brom_out <= 64'd7808447432725972242;
    12'd1395: brom_out <= 64'd829718688336966961;
    12'd883: brom_out <= 64'd2368990469369948360;
    12'd1907: brom_out <= 64'd7480559819299940365;
    12'd243: brom_out <= 64'd6012025652804998213;
    12'd1267: brom_out <= 64'd3008087335713497179;
    12'd755: brom_out <= 64'd8712593913693186332;
    12'd1779: brom_out <= 64'd2455840043548559201;
    12'd499: brom_out <= 64'd9049716330878161931;
    12'd1523: brom_out <= 64'd2880596291528857407;
    12'd1011: brom_out <= 64'd3481811138521427457;
    12'd2035: brom_out <= 64'd6478919389561179993;
    12'd11: brom_out <= 64'd5729530929914156035;
    12'd1035: brom_out <= 64'd6566468905650255250;
    12'd523: brom_out <= 64'd6385799882573814037;
    12'd1547: brom_out <= 64'd8910711434716434551;
    12'd267: brom_out <= 64'd4516276014168523495;
    12'd1291: brom_out <= 64'd145656868355011287;
    12'd779: brom_out <= 64'd4169901780951817161;
    12'd1803: brom_out <= 64'd905799661330999781;
    12'd139: brom_out <= 64'd4835634247680250719;
    12'd1163: brom_out <= 64'd6574981646075002534;
    12'd651: brom_out <= 64'd5584792192168107432;
    12'd1675: brom_out <= 64'd2752058282402856793;
    12'd395: brom_out <= 64'd8327204787394120192;
    12'd1419: brom_out <= 64'd5358308440264631809;
    12'd907: brom_out <= 64'd5893894784811767994;
    12'd1931: brom_out <= 64'd3942447305519050889;
    12'd75: brom_out <= 64'd8377901604773452116;
    12'd1099: brom_out <= 64'd6815651330881124184;
    12'd587: brom_out <= 64'd5227199790467636203;
    12'd1611: brom_out <= 64'd1509172337700286580;
    12'd331: brom_out <= 64'd7462029048422031806;
    12'd1355: brom_out <= 64'd8604485434315505735;
    12'd843: brom_out <= 64'd6414793489365941449;
    12'd1867: brom_out <= 64'd2393147964449530160;
    12'd203: brom_out <= 64'd7306856896100183088;
    12'd1227: brom_out <= 64'd4447745589333214354;
    12'd715: brom_out <= 64'd4498240959642217998;
    12'd1739: brom_out <= 64'd2058194682028382178;
    12'd459: brom_out <= 64'd1475031882489607674;
    12'd1483: brom_out <= 64'd4834804060714409564;
    12'd971: brom_out <= 64'd2538065853035112563;
    12'd1995: brom_out <= 64'd500197875907057540;
    12'd43: brom_out <= 64'd4918174515392184802;
    12'd1067: brom_out <= 64'd5776566466241365138;
    12'd555: brom_out <= 64'd680524271701586087;
    12'd1579: brom_out <= 64'd7926667544375359517;
    12'd299: brom_out <= 64'd790871527546262502;
    12'd1323: brom_out <= 64'd5421382544425298681;
    12'd811: brom_out <= 64'd1852964257181214603;
    12'd1835: brom_out <= 64'd1820466509108982119;
    12'd171: brom_out <= 64'd3577128854111046835;
    12'd1195: brom_out <= 64'd5932873316160418767;
    12'd683: brom_out <= 64'd2353401445000590928;
    12'd1707: brom_out <= 64'd694223862457378337;
    12'd427: brom_out <= 64'd360484740059425050;
    12'd1451: brom_out <= 64'd8228602517368847249;
    12'd939: brom_out <= 64'd3630606306430013653;
    12'd1963: brom_out <= 64'd2841349618467936928;
    12'd107: brom_out <= 64'd8641169949442141173;
    12'd1131: brom_out <= 64'd9178801026488190119;
    12'd619: brom_out <= 64'd6595457878857378400;
    12'd1643: brom_out <= 64'd3493839405849918059;
    12'd363: brom_out <= 64'd2850153989378393397;
    12'd1387: brom_out <= 64'd1460834046960258626;
    12'd875: brom_out <= 64'd2081215718459538783;
    12'd1899: brom_out <= 64'd3287110378832910730;
    12'd235: brom_out <= 64'd742784643922937883;
    12'd1259: brom_out <= 64'd8072235980992715391;
    12'd747: brom_out <= 64'd7909247277760472996;
    12'd1771: brom_out <= 64'd7389923767150689831;
    12'd491: brom_out <= 64'd4619850868153408086;
    12'd1515: brom_out <= 64'd2441840015076694878;
    12'd1003: brom_out <= 64'd6212407820719679929;
    12'd2027: brom_out <= 64'd7073835240576623789;
    12'd27: brom_out <= 64'd220500274699000058;
    12'd1051: brom_out <= 64'd3732354117739994962;
    12'd539: brom_out <= 64'd6421526328547564855;
    12'd1563: brom_out <= 64'd2530586432529640472;
    12'd283: brom_out <= 64'd4123312334176217225;
    12'd1307: brom_out <= 64'd9041130964638911268;
    12'd795: brom_out <= 64'd4566183379717796458;
    12'd1819: brom_out <= 64'd1757616478407663383;
    12'd155: brom_out <= 64'd2734242444567840901;
    12'd1179: brom_out <= 64'd3624582266943194900;
    12'd667: brom_out <= 64'd6786869815747781225;
    12'd1691: brom_out <= 64'd718743493023770566;
    12'd411: brom_out <= 64'd729810824920162793;
    12'd1435: brom_out <= 64'd1188276465581594610;
    12'd923: brom_out <= 64'd5139783655959744836;
    12'd1947: brom_out <= 64'd6900206609138170971;
    12'd91: brom_out <= 64'd1101597167942426836;
    12'd1115: brom_out <= 64'd605422831588364704;
    12'd603: brom_out <= 64'd4473474045233695924;
    12'd1627: brom_out <= 64'd5648624822793917853;
    12'd347: brom_out <= 64'd73717055544869389;
    12'd1371: brom_out <= 64'd1325625408625222270;
    12'd859: brom_out <= 64'd1776090422059416444;
    12'd1883: brom_out <= 64'd6819381790581932160;
    12'd219: brom_out <= 64'd2583420948749650888;
    12'd1243: brom_out <= 64'd1794510800470079672;
    12'd731: brom_out <= 64'd5102428610010320937;
    12'd1755: brom_out <= 64'd5223527647632959705;
    12'd475: brom_out <= 64'd3682180039723582694;
    12'd1499: brom_out <= 64'd8433275119812750687;
    12'd987: brom_out <= 64'd5112839996764513225;
    12'd2011: brom_out <= 64'd3856821850846535981;
    12'd59: brom_out <= 64'd3089285411360685289;
    12'd1083: brom_out <= 64'd2671675604543893083;
    12'd571: brom_out <= 64'd2290603348236949045;
    12'd1595: brom_out <= 64'd8727788904265190901;
    12'd315: brom_out <= 64'd6803294201327288707;
    12'd1339: brom_out <= 64'd1856831615331523383;
    12'd827: brom_out <= 64'd7770161374061953188;
    12'd1851: brom_out <= 64'd3256546726592676868;
    12'd187: brom_out <= 64'd7473753521031238993;
    12'd1211: brom_out <= 64'd8443274051820661742;
    12'd699: brom_out <= 64'd6688735190242104592;
    12'd1723: brom_out <= 64'd8595670644960839154;
    12'd443: brom_out <= 64'd7732607215987328911;
    12'd1467: brom_out <= 64'd8379321866420704450;
    12'd955: brom_out <= 64'd6945674550036316590;
    12'd1979: brom_out <= 64'd2535341830663400840;
    12'd123: brom_out <= 64'd5015573810118615339;
    12'd1147: brom_out <= 64'd8363836245864963634;
    12'd635: brom_out <= 64'd32125116951179213;
    12'd1659: brom_out <= 64'd7198242521742692345;
    12'd379: brom_out <= 64'd1235333264221809472;
    12'd1403: brom_out <= 64'd1928375831348488250;
    12'd891: brom_out <= 64'd8527425457839399944;
    12'd1915: brom_out <= 64'd6831933593153819906;
    12'd251: brom_out <= 64'd3545680560691756924;
    12'd1275: brom_out <= 64'd7718504265681008124;
    12'd763: brom_out <= 64'd7794858711406569316;
    12'd1787: brom_out <= 64'd6129983840930345678;
    12'd507: brom_out <= 64'd6969614548778718585;
    12'd1531: brom_out <= 64'd4846969929203527549;
    12'd1019: brom_out <= 64'd3023536135369317650;
    12'd2043: brom_out <= 64'd326945987357450470;
    12'd7: brom_out <= 64'd1196717673321766117;
    12'd1031: brom_out <= 64'd3491781143937178912;
    12'd519: brom_out <= 64'd4408752695654407648;
    12'd1543: brom_out <= 64'd5000700186948299879;
    12'd263: brom_out <= 64'd4219634770587921750;
    12'd1287: brom_out <= 64'd1320958211383417929;
    12'd775: brom_out <= 64'd682700647643264297;
    12'd1799: brom_out <= 64'd5444613374524628588;
    12'd135: brom_out <= 64'd1179502005020589858;
    12'd1159: brom_out <= 64'd6083514922364870232;
    12'd647: brom_out <= 64'd1809600597274552126;
    12'd1671: brom_out <= 64'd1024176671026003038;
    12'd391: brom_out <= 64'd4191546537857189221;
    12'd1415: brom_out <= 64'd2202724336846540116;
    12'd903: brom_out <= 64'd1877021610163541386;
    12'd1927: brom_out <= 64'd5995405915279804808;
    12'd71: brom_out <= 64'd6998202902482917701;
    12'd1095: brom_out <= 64'd1263511878798759381;
    12'd583: brom_out <= 64'd8021293061179377577;
    12'd1607: brom_out <= 64'd7582206566951821406;
    12'd327: brom_out <= 64'd4793887105630240660;
    12'd1351: brom_out <= 64'd1005982687865603721;
    12'd839: brom_out <= 64'd2183205339960394892;
    12'd1863: brom_out <= 64'd671045474484094746;
    12'd199: brom_out <= 64'd2464096157002094073;
    12'd1223: brom_out <= 64'd4698951168554923126;
    12'd711: brom_out <= 64'd5594102867212098478;
    12'd1735: brom_out <= 64'd3867060877188918314;
    12'd455: brom_out <= 64'd5729788999270214082;
    12'd1479: brom_out <= 64'd1029072485803360067;
    12'd967: brom_out <= 64'd3882434473969474706;
    12'd1991: brom_out <= 64'd6167912167594203538;
    12'd39: brom_out <= 64'd197803793147744096;
    12'd1063: brom_out <= 64'd3981789991754018619;
    12'd551: brom_out <= 64'd3513467328658626429;
    12'd1575: brom_out <= 64'd8525064474068460897;
    12'd295: brom_out <= 64'd3324554081399548856;
    12'd1319: brom_out <= 64'd946400147553460105;
    12'd807: brom_out <= 64'd3955913466213958211;
    12'd1831: brom_out <= 64'd1146971011575375733;
    12'd167: brom_out <= 64'd8758476752168223894;
    12'd1191: brom_out <= 64'd5016823419376867650;
    12'd679: brom_out <= 64'd6054674304173726790;
    12'd1703: brom_out <= 64'd4893994999723283549;
    12'd423: brom_out <= 64'd475642159627763285;
    12'd1447: brom_out <= 64'd7439733981079839283;
    12'd935: brom_out <= 64'd5543613125578900301;
    12'd1959: brom_out <= 64'd723257086799406522;
    12'd103: brom_out <= 64'd5580777950571297909;
    12'd1127: brom_out <= 64'd889628210544556757;
    12'd615: brom_out <= 64'd8209692884265780128;
    12'd1639: brom_out <= 64'd3168381531098261847;
    12'd359: brom_out <= 64'd1567032197242528000;
    12'd1383: brom_out <= 64'd8075643565788399825;
    12'd871: brom_out <= 64'd5576469314982004821;
    12'd1895: brom_out <= 64'd6212662201786385756;
    12'd231: brom_out <= 64'd1463997088774103234;
    12'd1255: brom_out <= 64'd5060595611919151390;
    12'd743: brom_out <= 64'd2151013669072265923;
    12'd1767: brom_out <= 64'd1854693964139895995;
    12'd487: brom_out <= 64'd7377995826428221440;
    12'd1511: brom_out <= 64'd7402617407341496296;
    12'd999: brom_out <= 64'd8799741510413925644;
    12'd2023: brom_out <= 64'd6684976454760300779;
    12'd23: brom_out <= 64'd8097826115473553654;
    12'd1047: brom_out <= 64'd1863936941917371814;
    12'd535: brom_out <= 64'd4070526297165743149;
    12'd1559: brom_out <= 64'd3699709539169764904;
    12'd279: brom_out <= 64'd8523351732208442783;
    12'd1303: brom_out <= 64'd4574373213825967675;
    12'd791: brom_out <= 64'd3625008606247825233;
    12'd1815: brom_out <= 64'd26440101996429966;
    12'd151: brom_out <= 64'd2269501464033279927;
    12'd1175: brom_out <= 64'd1077190625265622326;
    12'd663: brom_out <= 64'd1271420675811002564;
    12'd1687: brom_out <= 64'd7510039751267506069;
    12'd407: brom_out <= 64'd4059318855695747956;
    12'd1431: brom_out <= 64'd3347504886541291315;
    12'd919: brom_out <= 64'd7448472333334016475;
    12'd1943: brom_out <= 64'd1089436887455411285;
    12'd87: brom_out <= 64'd2555080649667943999;
    12'd1111: brom_out <= 64'd7066491535020407510;
    12'd599: brom_out <= 64'd8767220660621360094;
    12'd1623: brom_out <= 64'd8044165810467914666;
    12'd343: brom_out <= 64'd5797794430093649856;
    12'd1367: brom_out <= 64'd1335320839478398254;
    12'd855: brom_out <= 64'd372840657118470559;
    12'd1879: brom_out <= 64'd1290555543749468522;
    12'd215: brom_out <= 64'd5552602819486374918;
    12'd1239: brom_out <= 64'd7500467012641262154;
    12'd727: brom_out <= 64'd6521725718717934846;
    12'd1751: brom_out <= 64'd8681474579391462114;
    12'd471: brom_out <= 64'd8561448770356449495;
    12'd1495: brom_out <= 64'd2253915061275631925;
    12'd983: brom_out <= 64'd4472700481719007707;
    12'd2007: brom_out <= 64'd5771004432200253489;
    12'd55: brom_out <= 64'd4167850225838881549;
    12'd1079: brom_out <= 64'd1501599260911325108;
    12'd567: brom_out <= 64'd2431467625941313240;
    12'd1591: brom_out <= 64'd8557963212313699756;
    12'd311: brom_out <= 64'd9010706113524963170;
    12'd1335: brom_out <= 64'd6692702923211495212;
    12'd823: brom_out <= 64'd7981979497860488419;
    12'd1847: brom_out <= 64'd5970975953792141535;
    12'd183: brom_out <= 64'd8204676838312359150;
    12'd1207: brom_out <= 64'd1525782086824111198;
    12'd695: brom_out <= 64'd5983639989667179235;
    12'd1719: brom_out <= 64'd4661252615798978400;
    12'd439: brom_out <= 64'd7711398484518081392;
    12'd1463: brom_out <= 64'd2236578997351544867;
    12'd951: brom_out <= 64'd6924128837099585359;
    12'd1975: brom_out <= 64'd8963809510067359653;
    12'd119: brom_out <= 64'd5836581410912283100;
    12'd1143: brom_out <= 64'd7312806042340346359;
    12'd631: brom_out <= 64'd5002926744895353547;
    12'd1655: brom_out <= 64'd4907009643734143301;
    12'd375: brom_out <= 64'd5783583947165716781;
    12'd1399: brom_out <= 64'd7685848209204296144;
    12'd887: brom_out <= 64'd4403593538858485791;
    12'd1911: brom_out <= 64'd710478813732694724;
    12'd247: brom_out <= 64'd7063725616615073009;
    12'd1271: brom_out <= 64'd8846274975537736297;
    12'd759: brom_out <= 64'd7986402759624561996;
    12'd1783: brom_out <= 64'd6807047288131121316;
    12'd503: brom_out <= 64'd5592727481390712356;
    12'd1527: brom_out <= 64'd4364366340196051419;
    12'd1015: brom_out <= 64'd8797070563634888702;
    12'd2039: brom_out <= 64'd3000626997840900221;
    12'd15: brom_out <= 64'd2565707750441499058;
    12'd1039: brom_out <= 64'd7726711646517821485;
    12'd527: brom_out <= 64'd2996485441824910329;
    12'd1551: brom_out <= 64'd6256822282179377531;
    12'd271: brom_out <= 64'd8466905988399369262;
    12'd1295: brom_out <= 64'd6633789097031885863;
    12'd783: brom_out <= 64'd4429331098788724882;
    12'd1807: brom_out <= 64'd5432919712713374234;
    12'd143: brom_out <= 64'd6626098368862619876;
    12'd1167: brom_out <= 64'd2746605235690302343;
    12'd655: brom_out <= 64'd3742907819552853392;
    12'd1679: brom_out <= 64'd1457296783964949895;
    12'd399: brom_out <= 64'd2075815179298327183;
    12'd1423: brom_out <= 64'd4072091310264274448;
    12'd911: brom_out <= 64'd6013101536663769196;
    12'd1935: brom_out <= 64'd573479814256513508;
    12'd79: brom_out <= 64'd3622044979216983831;
    12'd1103: brom_out <= 64'd134034021807666817;
    12'd591: brom_out <= 64'd1127787708612535076;
    12'd1615: brom_out <= 64'd5423077958558031318;
    12'd335: brom_out <= 64'd8510449508983965512;
    12'd1359: brom_out <= 64'd1248384842966628456;
    12'd847: brom_out <= 64'd8792296984155581379;
    12'd1871: brom_out <= 64'd8373428133602290972;
    12'd207: brom_out <= 64'd1931047495115039244;
    12'd1231: brom_out <= 64'd5204721274885589650;
    12'd719: brom_out <= 64'd497959859408023041;
    12'd1743: brom_out <= 64'd4588670221998153173;
    12'd463: brom_out <= 64'd5265596843940117062;
    12'd1487: brom_out <= 64'd1160952030647706439;
    12'd975: brom_out <= 64'd3425575118838313248;
    12'd1999: brom_out <= 64'd2743982901281082008;
    12'd47: brom_out <= 64'd7361159851495798473;
    12'd1071: brom_out <= 64'd481102647340149789;
    12'd559: brom_out <= 64'd7231885404608803550;
    12'd1583: brom_out <= 64'd6438318227858851538;
    12'd303: brom_out <= 64'd2420540411133931766;
    12'd1327: brom_out <= 64'd1195686174748815171;
    12'd815: brom_out <= 64'd4065668864028310310;
    12'd1839: brom_out <= 64'd2362323282577995162;
    12'd175: brom_out <= 64'd4815692819958443175;
    12'd1199: brom_out <= 64'd3077747082406647727;
    12'd687: brom_out <= 64'd3828260745157223499;
    12'd1711: brom_out <= 64'd3986546580424101369;
    12'd431: brom_out <= 64'd3811253066581545128;
    12'd1455: brom_out <= 64'd7532977315832375559;
    12'd943: brom_out <= 64'd1665190001954023046;
    12'd1967: brom_out <= 64'd2098087234537064888;
    12'd111: brom_out <= 64'd828091323878167268;
    12'd1135: brom_out <= 64'd8544459384181573151;
    12'd623: brom_out <= 64'd5163228436461165095;
    12'd1647: brom_out <= 64'd6281474619484206548;
    12'd367: brom_out <= 64'd6990154071024195406;
    12'd1391: brom_out <= 64'd2937347601375647642;
    12'd879: brom_out <= 64'd7125465436638969639;
    12'd1903: brom_out <= 64'd7966166060157864076;
    12'd239: brom_out <= 64'd1119595535300504858;
    12'd1263: brom_out <= 64'd8164477216473543113;
    12'd751: brom_out <= 64'd4700788970051757419;
    12'd1775: brom_out <= 64'd6826850400113365008;
    12'd495: brom_out <= 64'd3952586212588864566;
    12'd1519: brom_out <= 64'd6450934739340643086;
    12'd1007: brom_out <= 64'd7605083119890874713;
    12'd2031: brom_out <= 64'd6848677136193455801;
    12'd31: brom_out <= 64'd4514273535597288556;
    12'd1055: brom_out <= 64'd5170043194338083281;
    12'd543: brom_out <= 64'd2535669803988329193;
    12'd1567: brom_out <= 64'd1609849005651730878;
    12'd287: brom_out <= 64'd3280335713029410903;
    12'd1311: brom_out <= 64'd6849064418324440089;
    12'd799: brom_out <= 64'd2828496737788716326;
    12'd1823: brom_out <= 64'd5844694662446046329;
    12'd159: brom_out <= 64'd2199597683219623913;
    12'd1183: brom_out <= 64'd7560298406862003465;
    12'd671: brom_out <= 64'd6885178931928983513;
    12'd1695: brom_out <= 64'd2531462407904144972;
    12'd415: brom_out <= 64'd5241450279032884119;
    12'd1439: brom_out <= 64'd4980098972437110768;
    12'd927: brom_out <= 64'd8064087142600323723;
    12'd1951: brom_out <= 64'd1288740745691906075;
    12'd95: brom_out <= 64'd4556586638489721473;
    12'd1119: brom_out <= 64'd1407137102196920649;
    12'd607: brom_out <= 64'd2513983781571577027;
    12'd1631: brom_out <= 64'd6371693099811397430;
    12'd351: brom_out <= 64'd2234213304222583316;
    12'd1375: brom_out <= 64'd7906729256064801356;
    12'd863: brom_out <= 64'd5074491527787452416;
    12'd1887: brom_out <= 64'd6718230231139610032;
    12'd223: brom_out <= 64'd1077895640556821346;
    12'd1247: brom_out <= 64'd8824798961944084459;
    12'd735: brom_out <= 64'd1959225301739326146;
    12'd1759: brom_out <= 64'd6001221512162512941;
    12'd479: brom_out <= 64'd8696952683898417962;
    12'd1503: brom_out <= 64'd6531887060912744218;
    12'd991: brom_out <= 64'd3521591547891566158;
    12'd2015: brom_out <= 64'd6146105024603525374;
    12'd63: brom_out <= 64'd7188693104123617185;
    12'd1087: brom_out <= 64'd3032780729918537940;
    12'd575: brom_out <= 64'd6094940225400254377;
    12'd1599: brom_out <= 64'd8564054125491362280;
    12'd319: brom_out <= 64'd7704680114262019375;
    12'd1343: brom_out <= 64'd8973803375737802424;
    12'd831: brom_out <= 64'd4461297653406609577;
    12'd1855: brom_out <= 64'd1716068777653910076;
    12'd191: brom_out <= 64'd6911963586344500087;
    12'd1215: brom_out <= 64'd6694492589769457580;
    12'd703: brom_out <= 64'd7325355971320287822;
    12'd1727: brom_out <= 64'd7060435521946386534;
    12'd447: brom_out <= 64'd81378846906711534;
    12'd1471: brom_out <= 64'd7931602618379434511;
    12'd959: brom_out <= 64'd8451356648349598988;
    12'd1983: brom_out <= 64'd6852251032093093684;
    12'd127: brom_out <= 64'd5015894486924318136;
    12'd1151: brom_out <= 64'd811675009939312370;
    12'd639: brom_out <= 64'd7188299900925906026;
    12'd1663: brom_out <= 64'd5460308741192036217;
    12'd383: brom_out <= 64'd3805511639449482562;
    12'd1407: brom_out <= 64'd2327897166772487923;
    12'd895: brom_out <= 64'd3443712695491297689;
    12'd1919: brom_out <= 64'd5922378199499929323;
    12'd255: brom_out <= 64'd8954848358245487830;
    12'd1279: brom_out <= 64'd27941890902324855;
    12'd767: brom_out <= 64'd6367475453121901558;
    12'd1791: brom_out <= 64'd3724189337875360527;
    12'd511: brom_out <= 64'd6363506754762091032;
    12'd1535: brom_out <= 64'd2280685463541578648;
    12'd1023: brom_out <= 64'd5743416372949675185;
    12'd2047: brom_out <= 64'd4423046145353804672;
    default: brom_out <= 64'h1;
    endcase
end

generate
    if(DELAY == 1) begin
        assign b = brom_out;
    end
endgenerate

endmodule

//-------------------------------------------------------------------------------------------------

module tw_rom_0_intt_nwc
#(
    parameter LOGN  = 0,
    parameter LOGQ  = 64,
    parameter DELAY = 1,
    parameter STAGE = 0
)(
    input            clk,
    input [LOGN-1:0] raddr,
    output[LOGQ-1:0] b
);

(* rom_style = "distributed" *)
reg [LOGQ-1:0] brom_out, brom_out2;

always @(posedge clk) begin
    case(raddr[0:0])
    1'd0: brom_out <= 64'd2672356941328551034;
    default: brom_out <= 64'h1;
    endcase
end

generate
    if(DELAY == 1) begin
        assign b = brom_out;
    end
endgenerate

endmodule

//-------------------------------------------------------------------------------------------------

module tw_rom_1_intt_nwc
#(
    parameter LOGN  = 1,
    parameter LOGQ  = 64,
    parameter DELAY = 1,
    parameter STAGE = 1
)(
    input            clk,
    input [LOGN-1:0] raddr,
    output[LOGQ-1:0] b
);

(* rom_style = "distributed" *)
reg [LOGQ-1:0] brom_out, brom_out2;

always @(posedge clk) begin
    case(raddr[STAGE-1:0])
    2'd0: brom_out <= 64'd5830754471805963540;
    2'd1: brom_out <= 64'd3247303257377812593;
    default: brom_out <= 64'h1;
    endcase
end

generate
    if(DELAY == 1) begin
        assign b = brom_out;
    end
endgenerate

endmodule

//-------------------------------------------------------------------------------------------------

module tw_rom_2_intt_nwc
#(
    parameter LOGN  = 2,
    parameter LOGQ  = 64,
    parameter DELAY = 1,
    parameter STAGE = 2
)(
    input            clk,
    input [LOGN-1:0] raddr,
    output[LOGQ-1:0] b
);

(* rom_style = "distributed" *)
reg [LOGQ-1:0] brom_out, brom_out2;

always @(posedge clk) begin
    case(raddr[STAGE-1:0])
    3'd0: brom_out <= 64'd8524270730790435434;
    3'd1: brom_out <= 64'd3430392906661205799;
    3'd2: brom_out <= 64'd6231927651766270000;
    3'd3: brom_out <= 64'd6341405124451893844;
    default: brom_out <= 64'h1;
    endcase
end

generate
    if(DELAY == 1) begin
        assign b = brom_out;
    end
endgenerate

endmodule

//-------------------------------------------------------------------------------------------------

module tw_rom_3_intt_nwc
#(
    parameter LOGN  = 3,
    parameter LOGQ  = 64,
    parameter DELAY = 1,
    parameter STAGE = 3
)(
    input            clk,
    input [LOGN-1:0] raddr,
    output[LOGQ-1:0] b
);

(* rom_style = "distributed" *)
reg [LOGQ-1:0] brom_out, brom_out2;

always @(posedge clk) begin
    case(raddr[STAGE-1:0])
    4'd0: brom_out <= 64'd7552580941491614922;
    4'd1: brom_out <= 64'd6420104328456603057;
    4'd2: brom_out <= 64'd1576457532180094608;
    4'd3: brom_out <= 64'd2075550771295400682;
    4'd4: brom_out <= 64'd8221312082853399401;
    4'd5: brom_out <= 64'd5156647865800837188;
    4'd6: brom_out <= 64'd3315193656759027728;
    4'd7: brom_out <= 64'd3306032853614922617;
    default: brom_out <= 64'h1;
    endcase
end

generate
    if(DELAY == 1) begin
        assign b = brom_out;
    end
endgenerate

endmodule

//-------------------------------------------------------------------------------------------------

module tw_rom_4_intt_nwc
#(
    parameter LOGN  = 4,
    parameter LOGQ  = 64,
    parameter DELAY = 1,
    parameter STAGE = 4
)(
    input            clk,
    input [LOGN-1:0] raddr,
    output[LOGQ-1:0] b
);

(* rom_style = "distributed" *)
reg [LOGQ-1:0] brom_out, brom_out2;

always @(posedge clk) begin
    case(raddr[STAGE-1:0])
    5'd0: brom_out <= 64'd8994868585466380386;
    5'd1: brom_out <= 64'd8158211732688145371;
    5'd2: brom_out <= 64'd4830110009435726389;
    5'd3: brom_out <= 64'd6179273730479935555;
    5'd4: brom_out <= 64'd37862187434532519;
    5'd5: brom_out <= 64'd6585485892914773929;
    5'd6: brom_out <= 64'd5675744442360421476;
    5'd7: brom_out <= 64'd5113008929590644365;
    5'd8: brom_out <= 64'd1299694352172497110;
    5'd9: brom_out <= 64'd6486214016837603816;
    5'd10: brom_out <= 64'd56701250192183654;
    5'd11: brom_out <= 64'd7598818098126613736;
    5'd12: brom_out <= 64'd4183627854902105294;
    5'd13: brom_out <= 64'd5349048256325193564;
    5'd14: brom_out <= 64'd350927547453619282;
    5'd15: brom_out <= 64'd517077598441490544;
    default: brom_out <= 64'h1;
    endcase
end

generate
    if(DELAY == 1) begin
        assign b = brom_out;
    end
endgenerate

endmodule

//-------------------------------------------------------------------------------------------------

module tw_rom_5_intt_nwc
#(
    parameter LOGN  = 5,
    parameter LOGQ  = 64,
    parameter DELAY = 1,
    parameter STAGE = 5
)(
    input            clk,
    input [LOGN-1:0] raddr,
    output[LOGQ-1:0] b
);

(* rom_style = "distributed" *)
reg [LOGQ-1:0] brom_out, brom_out2;

always @(posedge clk) begin
    case(raddr[STAGE-1:0])
    6'd0: brom_out <= 64'd8522641201658729225;
    6'd1: brom_out <= 64'd4312376496106318253;
    6'd2: brom_out <= 64'd3493420703660838670;
    6'd3: brom_out <= 64'd5700970638399166368;
    6'd4: brom_out <= 64'd220092981789821141;
    6'd5: brom_out <= 64'd4932371830946747484;
    6'd6: brom_out <= 64'd6754708753051563723;
    6'd7: brom_out <= 64'd7029009308789466914;
    6'd8: brom_out <= 64'd4096526975789124741;
    6'd9: brom_out <= 64'd3151400731738051651;
    6'd10: brom_out <= 64'd3568645759314256059;
    6'd11: brom_out <= 64'd3347897398381093651;
    6'd12: brom_out <= 64'd7594465691176760977;
    6'd13: brom_out <= 64'd8138265688407551998;
    6'd14: brom_out <= 64'd6553824577164106665;
    6'd15: brom_out <= 64'd3064886553006135361;
    6'd16: brom_out <= 64'd399907671399444804;
    6'd17: brom_out <= 64'd6219428817239726022;
    6'd18: brom_out <= 64'd7081664262943872385;
    6'd19: brom_out <= 64'd396810392799227093;
    6'd20: brom_out <= 64'd4387368684406258781;
    6'd21: brom_out <= 64'd913575703207508649;
    6'd22: brom_out <= 64'd7536036494695424491;
    6'd23: brom_out <= 64'd5272450513720306929;
    6'd24: brom_out <= 64'd9153529019070073013;
    6'd25: brom_out <= 64'd3627333257985458202;
    6'd26: brom_out <= 64'd1098418798196992532;
    6'd27: brom_out <= 64'd8487932953363879467;
    6'd28: brom_out <= 64'd9215155275265843933;
    6'd29: brom_out <= 64'd783439227444010058;
    6'd30: brom_out <= 64'd8939333164997474080;
    6'd31: brom_out <= 64'd2239006582231249492;
    default: brom_out <= 64'h1;
    endcase
end

generate
    if(DELAY == 1) begin
        assign b = brom_out;
    end
endgenerate

endmodule

//-------------------------------------------------------------------------------------------------

module tw_rom_6_intt_nwc
#(
    parameter LOGN  = 6,
    parameter LOGQ  = 64,
    parameter DELAY = 1,
    parameter STAGE = 6
)(
    input            clk,
    input [LOGN-1:0] raddr,
    output[LOGQ-1:0] b
);

(* rom_style = "distributed" *)
reg [LOGQ-1:0] brom_out, brom_out2;

always @(posedge clk) begin
    case(raddr[STAGE-1:0])
    7'd0: brom_out <= 64'd7109810547382757607;
    7'd1: brom_out <= 64'd367308847039914212;
    7'd2: brom_out <= 64'd7846670721510247656;
    7'd3: brom_out <= 64'd197869443449083407;
    7'd4: brom_out <= 64'd7395765625369856968;
    7'd5: brom_out <= 64'd2557533429584063773;
    7'd6: brom_out <= 64'd8045183738668174654;
    7'd7: brom_out <= 64'd2658841363941412644;
    7'd8: brom_out <= 64'd8427191891465618357;
    7'd9: brom_out <= 64'd5172951906572162055;
    7'd10: brom_out <= 64'd5664972945830873653;
    7'd11: brom_out <= 64'd3001368193782052215;
    7'd12: brom_out <= 64'd5695281814046274237;
    7'd13: brom_out <= 64'd7819862133573918962;
    7'd14: brom_out <= 64'd8684981881685669851;
    7'd15: brom_out <= 64'd1877889542523460400;
    7'd16: brom_out <= 64'd899388833242523160;
    7'd17: brom_out <= 64'd3203502557968907342;
    7'd18: brom_out <= 64'd2212575092587301459;
    7'd19: brom_out <= 64'd5696879247801395673;
    7'd20: brom_out <= 64'd2787040975931115558;
    7'd21: brom_out <= 64'd4781781563078534797;
    7'd22: brom_out <= 64'd4285083028815705402;
    7'd23: brom_out <= 64'd4649918672425962884;
    7'd24: brom_out <= 64'd1578301005375201442;
    7'd25: brom_out <= 64'd2765020618288638665;
    7'd26: brom_out <= 64'd3440773991301144844;
    7'd27: brom_out <= 64'd8678431911799834516;
    7'd28: brom_out <= 64'd1036407828749944283;
    7'd29: brom_out <= 64'd186723147937826347;
    7'd30: brom_out <= 64'd6694132473816219222;
    7'd31: brom_out <= 64'd3569994870397592703;
    7'd32: brom_out <= 64'd2221241477869573467;
    7'd33: brom_out <= 64'd5624992943020008915;
    7'd34: brom_out <= 64'd4303776052874420108;
    7'd35: brom_out <= 64'd9002203609698631477;
    7'd36: brom_out <= 64'd1227696580085511339;
    7'd37: brom_out <= 64'd2136919832022164317;
    7'd38: brom_out <= 64'd3278507459918854810;
    7'd39: brom_out <= 64'd1153068650459044761;
    7'd40: brom_out <= 64'd8848016001656751714;
    7'd41: brom_out <= 64'd7006916387714091417;
    7'd42: brom_out <= 64'd6107523945568620274;
    7'd43: brom_out <= 64'd6297296671813620711;
    7'd44: brom_out <= 64'd3751399568142705465;
    7'd45: brom_out <= 64'd4860367702623205232;
    7'd46: brom_out <= 64'd6519545547382872352;
    7'd47: brom_out <= 64'd2597310436694665440;
    7'd48: brom_out <= 64'd5942845905398696661;
    7'd49: brom_out <= 64'd5139493591777994574;
    7'd50: brom_out <= 64'd7668063874127122800;
    7'd51: brom_out <= 64'd4505979271650606453;
    7'd52: brom_out <= 64'd8916215354504105080;
    7'd53: brom_out <= 64'd4512407425411054796;
    7'd54: brom_out <= 64'd146455696100183948;
    7'd55: brom_out <= 64'd1049049003178351694;
    7'd56: brom_out <= 64'd3330099465632933800;
    7'd57: brom_out <= 64'd3904396817663497520;
    7'd58: brom_out <= 64'd2941708752279192580;
    7'd59: brom_out <= 64'd8004307236827214629;
    7'd60: brom_out <= 64'd6960102488200083335;
    7'd61: brom_out <= 64'd7951696391921209588;
    7'd62: brom_out <= 64'd5182472792701730007;
    7'd63: brom_out <= 64'd8953373582369623737;
    default: brom_out <= 64'h1;
    endcase
end

generate
    if(DELAY == 1) begin
        assign b = brom_out;
    end
endgenerate

endmodule

//-------------------------------------------------------------------------------------------------

module tw_rom_7_intt_nwc
#(
    parameter LOGN  = 7,
    parameter LOGQ  = 64,
    parameter DELAY = 1,
    parameter STAGE = 7
)(
    input            clk,
    input [LOGN-1:0] raddr,
    output[LOGQ-1:0] b
);

(* rom_style = "distributed" *)
reg [LOGQ-1:0] brom_out, brom_out2;

always @(posedge clk) begin
    case(raddr[STAGE-1:0])
    8'd0: brom_out <= 64'd1954326138506476951;
    8'd1: brom_out <= 64'd4331403685672425430;
    8'd2: brom_out <= 64'd3283704730850768061;
    8'd3: brom_out <= 64'd4689801662437794854;
    8'd4: brom_out <= 64'd1550373778486368231;
    8'd5: brom_out <= 64'd5152867596778053751;
    8'd6: brom_out <= 64'd3350265901562279742;
    8'd7: brom_out <= 64'd7316289197091491357;
    8'd8: brom_out <= 64'd5103863865215982985;
    8'd9: brom_out <= 64'd3979599900047654998;
    8'd10: brom_out <= 64'd4459335126207999102;
    8'd11: brom_out <= 64'd8606842531585174143;
    8'd12: brom_out <= 64'd425055851346828692;
    8'd13: brom_out <= 64'd4604048451863389211;
    8'd14: brom_out <= 64'd5144400845762011825;
    8'd15: brom_out <= 64'd1186334652025577480;
    8'd16: brom_out <= 64'd3800020316465466232;
    8'd17: brom_out <= 64'd3477229189222177394;
    8'd18: brom_out <= 64'd530820408317780081;
    8'd19: brom_out <= 64'd3911674197792430825;
    8'd20: brom_out <= 64'd7581449063832142145;
    8'd21: brom_out <= 64'd2515433623371240219;
    8'd22: brom_out <= 64'd2648394196747926594;
    8'd23: brom_out <= 64'd5856315971097697291;
    8'd24: brom_out <= 64'd4049949528056965473;
    8'd25: brom_out <= 64'd3929914254541433141;
    8'd26: brom_out <= 64'd3232312203174602576;
    8'd27: brom_out <= 64'd7377924364550459486;
    8'd28: brom_out <= 64'd2373934992687024350;
    8'd29: brom_out <= 64'd8484153087462644695;
    8'd30: brom_out <= 64'd116462860189362305;
    8'd31: brom_out <= 64'd308674020057320967;
    8'd32: brom_out <= 64'd1751956540902519909;
    8'd33: brom_out <= 64'd4555648174004762903;
    8'd34: brom_out <= 64'd4303621306168106290;
    8'd35: brom_out <= 64'd3777108908419357151;
    8'd36: brom_out <= 64'd4373689981798860983;
    8'd37: brom_out <= 64'd5850377550468370218;
    8'd38: brom_out <= 64'd8538732393051528922;
    8'd39: brom_out <= 64'd3540997547282744152;
    8'd40: brom_out <= 64'd8711844274856048743;
    8'd41: brom_out <= 64'd7767534610063544800;
    8'd42: brom_out <= 64'd8473011002040519090;
    8'd43: brom_out <= 64'd3511217556398212621;
    8'd44: brom_out <= 64'd2597193474166918635;
    8'd45: brom_out <= 64'd1294300835907513996;
    8'd46: brom_out <= 64'd7270528764703572049;
    8'd47: brom_out <= 64'd2848104795771373212;
    8'd48: brom_out <= 64'd5608244685349795074;
    8'd49: brom_out <= 64'd1481448112490312089;
    8'd50: brom_out <= 64'd2673146875957441753;
    8'd51: brom_out <= 64'd4911251316354890590;
    8'd52: brom_out <= 64'd6115453565595858482;
    8'd53: brom_out <= 64'd2394991428284228318;
    8'd54: brom_out <= 64'd4182528396652029681;
    8'd55: brom_out <= 64'd6904336388986369203;
    8'd56: brom_out <= 64'd4783446724181950094;
    8'd57: brom_out <= 64'd4222427797676162143;
    8'd58: brom_out <= 64'd525772590065176804;
    8'd59: brom_out <= 64'd7357982398955724706;
    8'd60: brom_out <= 64'd2240676235245539362;
    8'd61: brom_out <= 64'd8045933869221030274;
    8'd62: brom_out <= 64'd3540330357633574851;
    8'd63: brom_out <= 64'd189984415773888079;
    8'd64: brom_out <= 64'd638376895518254818;
    8'd65: brom_out <= 64'd213963717958513684;
    8'd66: brom_out <= 64'd6983082545545823820;
    8'd67: brom_out <= 64'd1475184694732677003;
    8'd68: brom_out <= 64'd8353545677674474114;
    8'd69: brom_out <= 64'd7990717558823176439;
    8'd70: brom_out <= 64'd7385691322947166451;
    8'd71: brom_out <= 64'd8983301363007214294;
    8'd72: brom_out <= 64'd61021348019496634;
    8'd73: brom_out <= 64'd7199727630968781876;
    8'd74: brom_out <= 64'd4014557695810220726;
    8'd75: brom_out <= 64'd1934046995492470519;
    8'd76: brom_out <= 64'd1517542463022799200;
    8'd77: brom_out <= 64'd8413885842224603145;
    8'd78: brom_out <= 64'd877801006820804151;
    8'd79: brom_out <= 64'd6414683792461298086;
    8'd80: brom_out <= 64'd4219842663924998847;
    8'd81: brom_out <= 64'd6420309666027690116;
    8'd82: brom_out <= 64'd3804932470683584806;
    8'd83: brom_out <= 64'd9216323394984268281;
    8'd84: brom_out <= 64'd6299957421132029054;
    8'd85: brom_out <= 64'd3539296286503267835;
    8'd86: brom_out <= 64'd404908965326887961;
    8'd87: brom_out <= 64'd5691952397696844857;
    8'd88: brom_out <= 64'd998199631558019834;
    8'd89: brom_out <= 64'd5858083699088023850;
    8'd90: brom_out <= 64'd4598077949735866368;
    8'd91: brom_out <= 64'd4286709743008445481;
    8'd92: brom_out <= 64'd2298000442561295564;
    8'd93: brom_out <= 64'd53012713845076886;
    8'd94: brom_out <= 64'd6668987832474222721;
    8'd95: brom_out <= 64'd8413311218309265442;
    8'd96: brom_out <= 64'd8724403251150692469;
    8'd97: brom_out <= 64'd1072204180962969925;
    8'd98: brom_out <= 64'd5063682243788939407;
    8'd99: brom_out <= 64'd1282785490896801108;
    8'd100: brom_out <= 64'd7676640257482938795;
    8'd101: brom_out <= 64'd3902463277252418616;
    8'd102: brom_out <= 64'd9165811856331148261;
    8'd103: brom_out <= 64'd3989946030105363693;
    8'd104: brom_out <= 64'd7083682629857346686;
    8'd105: brom_out <= 64'd3616208387143208215;
    8'd106: brom_out <= 64'd2049717196365692321;
    8'd107: brom_out <= 64'd5636376557987066388;
    8'd108: brom_out <= 64'd6159062186366994793;
    8'd109: brom_out <= 64'd3504504943674790294;
    8'd110: brom_out <= 64'd4610082520291612538;
    8'd111: brom_out <= 64'd7238891700725414957;
    8'd112: brom_out <= 64'd3233457307195839204;
    8'd113: brom_out <= 64'd7605304680211549935;
    8'd114: brom_out <= 64'd6157433478933926008;
    8'd115: brom_out <= 64'd6074144695585879373;
    8'd116: brom_out <= 64'd7732484480248053853;
    8'd117: brom_out <= 64'd5620168497870933020;
    8'd118: brom_out <= 64'd4540514741108745753;
    8'd119: brom_out <= 64'd5662252708010606551;
    8'd120: brom_out <= 64'd1003412244194710405;
    8'd121: brom_out <= 64'd9000403498996357728;
    8'd122: brom_out <= 64'd8100974381305375741;
    8'd123: brom_out <= 64'd370750906239421062;
    8'd124: brom_out <= 64'd1744224572002386106;
    8'd125: brom_out <= 64'd8630329754039042439;
    8'd126: brom_out <= 64'd5426989541722031372;
    8'd127: brom_out <= 64'd7923915991122322492;
    default: brom_out <= 64'h1;
    endcase
end

generate
    if(DELAY == 1) begin
        assign b = brom_out;
    end
endgenerate

endmodule

//-------------------------------------------------------------------------------------------------

module tw_rom_8_intt_nwc
#(
    parameter LOGN  = 8,
    parameter LOGQ  = 64,
    parameter DELAY = 1,
    parameter STAGE = 8
)(
    input            clk,
    input [LOGN-1:0] raddr,
    output[LOGQ-1:0] b
);

(* ram_style = "block" *)
reg [LOGQ-1:0] brom_out, brom_out2;

always @(posedge clk) begin
    case(raddr[STAGE-1:0])
    9'd0: brom_out <= 64'd589261252211951087;
    9'd1: brom_out <= 64'd4077894327936387370;
    9'd2: brom_out <= 64'd6288258031243589040;
    9'd3: brom_out <= 64'd6308906059119793794;
    9'd4: brom_out <= 64'd1692640787285258321;
    9'd5: brom_out <= 64'd1619821793978715171;
    9'd6: brom_out <= 64'd419593050970393370;
    9'd7: brom_out <= 64'd6191527649035338270;
    9'd8: brom_out <= 64'd4699798339353139954;
    9'd9: brom_out <= 64'd6908457582704881495;
    9'd10: brom_out <= 64'd25503325735103202;
    9'd11: brom_out <= 64'd4687870931622476041;
    9'd12: brom_out <= 64'd3069294723345492836;
    9'd13: brom_out <= 64'd2808246389382168329;
    9'd14: brom_out <= 64'd4640137479215230119;
    9'd15: brom_out <= 64'd118759412684387883;
    9'd16: brom_out <= 64'd3815069067454082137;
    9'd17: brom_out <= 64'd6092909804324845418;
    9'd18: brom_out <= 64'd4399302856811857180;
    9'd19: brom_out <= 64'd2213917089242083356;
    9'd20: brom_out <= 64'd4541598978652527422;
    9'd21: brom_out <= 64'd1146302675032785038;
    9'd22: brom_out <= 64'd8402264118125672286;
    9'd23: brom_out <= 64'd5339911404069392687;
    9'd24: brom_out <= 64'd6623073124285805253;
    9'd25: brom_out <= 64'd6871996863026178947;
    9'd26: brom_out <= 64'd1123077664257713665;
    9'd27: brom_out <= 64'd7040469710198952938;
    9'd28: brom_out <= 64'd778504295643026436;
    9'd29: brom_out <= 64'd1967349882660717137;
    9'd30: brom_out <= 64'd9112039889942036181;
    9'd31: brom_out <= 64'd3443976834896946719;
    9'd32: brom_out <= 64'd105711516313429415;
    9'd33: brom_out <= 64'd103409383105209966;
    9'd34: brom_out <= 64'd4809545509471822219;
    9'd35: brom_out <= 64'd3921481593659637310;
    9'd36: brom_out <= 64'd63319580882334172;
    9'd37: brom_out <= 64'd6201111492212702581;
    9'd38: brom_out <= 64'd5883112818552593198;
    9'd39: brom_out <= 64'd9050257226618106939;
    9'd40: brom_out <= 64'd3810478311941277648;
    9'd41: brom_out <= 64'd7522099694907264830;
    9'd42: brom_out <= 64'd5631173395608091303;
    9'd43: brom_out <= 64'd5744306578764950661;
    9'd44: brom_out <= 64'd13835922099275263;
    9'd45: brom_out <= 64'd6560069435788688786;
    9'd46: brom_out <= 64'd2119102014119758127;
    9'd47: brom_out <= 64'd8431074821866737843;
    9'd48: brom_out <= 64'd3074762226706504168;
    9'd49: brom_out <= 64'd7007767720959207427;
    9'd50: brom_out <= 64'd3733077519005931989;
    9'd51: brom_out <= 64'd8474334919647044364;
    9'd52: brom_out <= 64'd2762686794518083477;
    9'd53: brom_out <= 64'd1095734946061864758;
    9'd54: brom_out <= 64'd4717167128727700595;
    9'd55: brom_out <= 64'd3322932605445341239;
    9'd56: brom_out <= 64'd4424637403257552821;
    9'd57: brom_out <= 64'd8163823191960297400;
    9'd58: brom_out <= 64'd8988229203291965646;
    9'd59: brom_out <= 64'd1300031822741507656;
    9'd60: brom_out <= 64'd3154929291392879223;
    9'd61: brom_out <= 64'd2319697542307896639;
    9'd62: brom_out <= 64'd514747083188271512;
    9'd63: brom_out <= 64'd4457485840176994766;
    9'd64: brom_out <= 64'd2304407482455379602;
    9'd65: brom_out <= 64'd4039054657987158917;
    9'd66: brom_out <= 64'd7050015494578529162;
    9'd67: brom_out <= 64'd5036136080121317251;
    9'd68: brom_out <= 64'd2593142759304359169;
    9'd69: brom_out <= 64'd2123928139285501187;
    9'd70: brom_out <= 64'd7186780195665525402;
    9'd71: brom_out <= 64'd7795526000590093317;
    9'd72: brom_out <= 64'd8381422672956537638;
    9'd73: brom_out <= 64'd2826957597084985722;
    9'd74: brom_out <= 64'd3672256128084492157;
    9'd75: brom_out <= 64'd7438283622837626809;
    9'd76: brom_out <= 64'd4289143564906162427;
    9'd77: brom_out <= 64'd3043838015584556076;
    9'd78: brom_out <= 64'd3205821663686069884;
    9'd79: brom_out <= 64'd1320831224533501879;
    9'd80: brom_out <= 64'd5859805713605662769;
    9'd81: brom_out <= 64'd1522999986540185734;
    9'd82: brom_out <= 64'd4973940462469037197;
    9'd83: brom_out <= 64'd6205769828923989477;
    9'd84: brom_out <= 64'd1196742974566397564;
    9'd85: brom_out <= 64'd2755115531749018871;
    9'd86: brom_out <= 64'd1938893570832931913;
    9'd87: brom_out <= 64'd2925505979841076067;
    9'd88: brom_out <= 64'd8246503946328159541;
    9'd89: brom_out <= 64'd3330517986526407221;
    9'd90: brom_out <= 64'd9147405191682765924;
    9'd91: brom_out <= 64'd3533540111080492141;
    9'd92: brom_out <= 64'd7655235938190610575;
    9'd93: brom_out <= 64'd4428743309412020209;
    9'd94: brom_out <= 64'd2760205288818577340;
    9'd95: brom_out <= 64'd642165299275900477;
    9'd96: brom_out <= 64'd6140091155236073342;
    9'd97: brom_out <= 64'd4246734587113910045;
    9'd98: brom_out <= 64'd8568619109861133075;
    9'd99: brom_out <= 64'd334488714186208727;
    9'd100: brom_out <= 64'd7432579756332737374;
    9'd101: brom_out <= 64'd3000563892240665083;
    9'd102: brom_out <= 64'd1391934389550943589;
    9'd103: brom_out <= 64'd2097737965174890192;
    9'd104: brom_out <= 64'd5493607054285716978;
    9'd105: brom_out <= 64'd2994197068779524467;
    9'd106: brom_out <= 64'd7276128854935879606;
    9'd107: brom_out <= 64'd7166058291707821460;
    9'd108: brom_out <= 64'd8831854030073042443;
    9'd109: brom_out <= 64'd789883360842779651;
    9'd110: brom_out <= 64'd2390447308213969615;
    9'd111: brom_out <= 64'd2071065103091007619;
    9'd112: brom_out <= 64'd724665762548809205;
    9'd113: brom_out <= 64'd6438983336492458386;
    9'd114: brom_out <= 64'd6479075097794724567;
    9'd115: brom_out <= 64'd8318711696260686832;
    9'd116: brom_out <= 64'd2118560143660212305;
    9'd117: brom_out <= 64'd1181817984886545321;
    9'd118: brom_out <= 64'd288492233688630408;
    9'd119: brom_out <= 64'd6314487893858783218;
    9'd120: brom_out <= 64'd679541861932208943;
    9'd121: brom_out <= 64'd2573214998270751675;
    9'd122: brom_out <= 64'd6696074260904623189;
    9'd123: brom_out <= 64'd8952875239077973570;
    9'd124: brom_out <= 64'd1685264228382100567;
    9'd125: brom_out <= 64'd4042041304395522620;
    9'd126: brom_out <= 64'd9208128174980151621;
    9'd127: brom_out <= 64'd1009423597135954028;
    9'd128: brom_out <= 64'd5387988075752117001;
    9'd129: brom_out <= 64'd3633169461159069704;
    9'd130: brom_out <= 64'd6055615886165633566;
    9'd131: brom_out <= 64'd7478733514354970269;
    9'd132: brom_out <= 64'd2274224641090761133;
    9'd133: brom_out <= 64'd7926032648594701020;
    9'd134: brom_out <= 64'd6112812087681150717;
    9'd135: brom_out <= 64'd6125288382695497236;
    9'd136: brom_out <= 64'd2342259468597363952;
    9'd137: brom_out <= 64'd1245574904084707370;
    9'd138: brom_out <= 64'd7731827774365937206;
    9'd139: brom_out <= 64'd7232379796619682380;
    9'd140: brom_out <= 64'd7964702205624645653;
    9'd141: brom_out <= 64'd5712954573871062153;
    9'd142: brom_out <= 64'd7764378251476652588;
    9'd143: brom_out <= 64'd8923477083739365998;
    9'd144: brom_out <= 64'd5482795640382241052;
    9'd145: brom_out <= 64'd2461761240587664975;
    9'd146: brom_out <= 64'd2087675356032182493;
    9'd147: brom_out <= 64'd8734263905964823460;
    9'd148: brom_out <= 64'd2489664880988935793;
    9'd149: brom_out <= 64'd588990440229857487;
    9'd150: brom_out <= 64'd5534417286816936371;
    9'd151: brom_out <= 64'd7936222448925179441;
    9'd152: brom_out <= 64'd4083084011917672932;
    9'd153: brom_out <= 64'd4767163061551348798;
    9'd154: brom_out <= 64'd1353263455556178614;
    9'd155: brom_out <= 64'd7925835341717889611;
    9'd156: brom_out <= 64'd7546502125228201480;
    9'd157: brom_out <= 64'd8229307188733692697;
    9'd158: brom_out <= 64'd5375797780357178476;
    9'd159: brom_out <= 64'd6923531029202165725;
    9'd160: brom_out <= 64'd6206391997638971135;
    9'd161: brom_out <= 64'd5563390978648112997;
    9'd162: brom_out <= 64'd6406968088848326056;
    9'd163: brom_out <= 64'd2268769362602750940;
    9'd164: brom_out <= 64'd9025136229324579910;
    9'd165: brom_out <= 64'd3528013818440306228;
    9'd166: brom_out <= 64'd4144380039276126840;
    9'd167: brom_out <= 64'd4876670574342399508;
    9'd168: brom_out <= 64'd4261452167139972416;
    9'd169: brom_out <= 64'd7908385913244527825;
    9'd170: brom_out <= 64'd3996836862911863169;
    9'd171: brom_out <= 64'd1229607629888877110;
    9'd172: brom_out <= 64'd828204405032100156;
    9'd173: brom_out <= 64'd8201782537523154361;
    9'd174: brom_out <= 64'd5995689611450984939;
    9'd175: brom_out <= 64'd4890576512707660646;
    9'd176: brom_out <= 64'd8341990074231113286;
    9'd177: brom_out <= 64'd2886148160064218946;
    9'd178: brom_out <= 64'd9003283877010505837;
    9'd179: brom_out <= 64'd4864032996040264162;
    9'd180: brom_out <= 64'd493093305913360701;
    9'd181: brom_out <= 64'd6104570640463597240;
    9'd182: brom_out <= 64'd4198473183879260811;
    9'd183: brom_out <= 64'd2069829275119115364;
    9'd184: brom_out <= 64'd7207482519161478029;
    9'd185: brom_out <= 64'd5112830294521799360;
    9'd186: brom_out <= 64'd1689880283676574380;
    9'd187: brom_out <= 64'd8679794296778572036;
    9'd188: brom_out <= 64'd2424707082823665464;
    9'd189: brom_out <= 64'd1209549302495265994;
    9'd190: brom_out <= 64'd6983160120422035266;
    9'd191: brom_out <= 64'd1289000951569658236;
    9'd192: brom_out <= 64'd2136168651708792999;
    9'd193: brom_out <= 64'd2790823145095613708;
    9'd194: brom_out <= 64'd480039465659720163;
    9'd195: brom_out <= 64'd2237522202805299556;
    9'd196: brom_out <= 64'd4211385562664614622;
    9'd197: brom_out <= 64'd1403394617657524198;
    9'd198: brom_out <= 64'd3424547160011928515;
    9'd199: brom_out <= 64'd8821413667448041115;
    9'd200: brom_out <= 64'd3042305502217840860;
    9'd201: brom_out <= 64'd1114624846972672018;
    9'd202: brom_out <= 64'd4713107804338707145;
    9'd203: brom_out <= 64'd2674968781932012466;
    9'd204: brom_out <= 64'd4854671826706628546;
    9'd205: brom_out <= 64'd8370295069151698855;
    9'd206: brom_out <= 64'd4638332250641664029;
    9'd207: brom_out <= 64'd7257217136825855779;
    9'd208: brom_out <= 64'd4084274140532747064;
    9'd209: brom_out <= 64'd7840499756043601545;
    9'd210: brom_out <= 64'd1630151818050992230;
    9'd211: brom_out <= 64'd3070088855073214330;
    9'd212: brom_out <= 64'd1172075295808189902;
    9'd213: brom_out <= 64'd1282831678063137055;
    9'd214: brom_out <= 64'd2369054697196546747;
    9'd215: brom_out <= 64'd7060379826744834670;
    9'd216: brom_out <= 64'd975391933298444430;
    9'd217: brom_out <= 64'd1419718399260074455;
    9'd218: brom_out <= 64'd3414595762090462243;
    9'd219: brom_out <= 64'd3867037900001858642;
    9'd220: brom_out <= 64'd120958337512701340;
    9'd221: brom_out <= 64'd431852270420361886;
    9'd222: brom_out <= 64'd2126423270618795487;
    9'd223: brom_out <= 64'd7100305522130918214;
    9'd224: brom_out <= 64'd2309488133539518628;
    9'd225: brom_out <= 64'd2269490171363922800;
    9'd226: brom_out <= 64'd329757546751791319;
    9'd227: brom_out <= 64'd8255979094666319636;
    9'd228: brom_out <= 64'd2992419980413818290;
    9'd229: brom_out <= 64'd5090820233960942835;
    9'd230: brom_out <= 64'd7674084484962021186;
    9'd231: brom_out <= 64'd3673423285967211399;
    9'd232: brom_out <= 64'd6947418755193653346;
    9'd233: brom_out <= 64'd6735392153401256686;
    9'd234: brom_out <= 64'd2139948861091713406;
    9'd235: brom_out <= 64'd6211254294135545461;
    9'd236: brom_out <= 64'd5754639100736438191;
    9'd237: brom_out <= 64'd2295357414439001689;
    9'd238: brom_out <= 64'd6880027384668613344;
    9'd239: brom_out <= 64'd6713575814653797923;
    9'd240: brom_out <= 64'd2954926496463500137;
    9'd241: brom_out <= 64'd846427375569667325;
    9'd242: brom_out <= 64'd3509794690809297077;
    9'd243: brom_out <= 64'd7624377972788189806;
    9'd244: brom_out <= 64'd6465598422296266431;
    9'd245: brom_out <= 64'd7611478067078673454;
    9'd246: brom_out <= 64'd1229558861263779893;
    9'd247: brom_out <= 64'd4831330309061259958;
    9'd248: brom_out <= 64'd8568248147423400136;
    9'd249: brom_out <= 64'd4771080522426822960;
    9'd250: brom_out <= 64'd5040072808927960902;
    9'd251: brom_out <= 64'd6297962505593583257;
    9'd252: brom_out <= 64'd6993322709341685228;
    9'd253: brom_out <= 64'd3161501911437101950;
    9'd254: brom_out <= 64'd571056314985110660;
    9'd255: brom_out <= 64'd1617878164001618876;
    default: brom_out <= 64'h1;
    endcase
end

generate
    if(DELAY == 1) begin
        assign b = brom_out;
    end
endgenerate

endmodule

//-------------------------------------------------------------------------------------------------

module tw_rom_9_intt_nwc
#(
    parameter LOGN  = 9,
    parameter LOGQ  = 64,
    parameter DELAY = 1,
    parameter STAGE = 9
)(
    input            clk,
    input [LOGN-1:0] raddr,
    output[LOGQ-1:0] b
);

(* ram_style = "block" *)
reg [LOGQ-1:0] brom_out, brom_out2;

always @(posedge clk) begin
    case(raddr[STAGE-1:0])
    10'd0: brom_out <= 64'd4419823402085286805;
    10'd1: brom_out <= 64'd1302461877294294752;
    10'd2: brom_out <= 64'd1530441695513114145;
    10'd3: brom_out <= 64'd1148748572447853663;
    10'd4: brom_out <= 64'd591599354290729504;
    10'd5: brom_out <= 64'd2128688671372429517;
    10'd6: brom_out <= 64'd2637825524469816123;
    10'd7: brom_out <= 64'd7827055078403768749;
    10'd8: brom_out <= 64'd126780732691162523;
    10'd9: brom_out <= 64'd8422066526749857360;
    10'd10: brom_out <= 64'd2453400897160557404;
    10'd11: brom_out <= 64'd6930291399587126145;
    10'd12: brom_out <= 64'd4267549409682314842;
    10'd13: brom_out <= 64'd2564632701129035616;
    10'd14: brom_out <= 64'd2841282234719890953;
    10'd15: brom_out <= 64'd7675678812830399463;
    10'd16: brom_out <= 64'd1375366390208185636;
    10'd17: brom_out <= 64'd2333492359452369891;
    10'd18: brom_out <= 64'd8081529454545222189;
    10'd19: brom_out <= 64'd7501208786978008007;
    10'd20: brom_out <= 64'd5819278190607705101;
    10'd21: brom_out <= 64'd2303593298178961587;
    10'd22: brom_out <= 64'd6474362064501644335;
    10'd23: brom_out <= 64'd4736437786329405404;
    10'd24: brom_out <= 64'd2506455365048153705;
    10'd25: brom_out <= 64'd464207075437736585;
    10'd26: brom_out <= 64'd5718898105580234973;
    10'd27: brom_out <= 64'd1525969772597555080;
    10'd28: brom_out <= 64'd71856063203078695;
    10'd29: brom_out <= 64'd6758808554109629452;
    10'd30: brom_out <= 64'd8374065344585748418;
    10'd31: brom_out <= 64'd513197978269968746;
    10'd32: brom_out <= 64'd8890008476498274928;
    10'd33: brom_out <= 64'd9055069812194889269;
    10'd34: brom_out <= 64'd2192817591669103432;
    10'd35: brom_out <= 64'd8100239580842297638;
    10'd36: brom_out <= 64'd2812120985173393103;
    10'd37: brom_out <= 64'd2869653304992504690;
    10'd38: brom_out <= 64'd5631842603051479664;
    10'd39: brom_out <= 64'd3909124456639709257;
    10'd40: brom_out <= 64'd4191157764168893931;
    10'd41: brom_out <= 64'd8054775185533533641;
    10'd42: brom_out <= 64'd5789862131438988414;
    10'd43: brom_out <= 64'd7638000315786716856;
    10'd44: brom_out <= 64'd275704973706589048;
    10'd45: brom_out <= 64'd3188911167348901112;
    10'd46: brom_out <= 64'd8411137007651424480;
    10'd47: brom_out <= 64'd2164694949571207915;
    10'd48: brom_out <= 64'd8623641753162776723;
    10'd49: brom_out <= 64'd6614846501772335324;
    10'd50: brom_out <= 64'd3023699520674774026;
    10'd51: brom_out <= 64'd1202062708655863367;
    10'd52: brom_out <= 64'd3772604775828423211;
    10'd53: brom_out <= 64'd4809087518643142365;
    10'd54: brom_out <= 64'd4400563506437680864;
    10'd55: brom_out <= 64'd279308063968193427;
    10'd56: brom_out <= 64'd2441744474732892698;
    10'd57: brom_out <= 64'd3864252773300489849;
    10'd58: brom_out <= 64'd8144458466683990449;
    10'd59: brom_out <= 64'd4400937907073847735;
    10'd60: brom_out <= 64'd6994819051443280820;
    10'd61: brom_out <= 64'd3821757200135596825;
    10'd62: brom_out <= 64'd1388160391904732628;
    10'd63: brom_out <= 64'd4110788945313777124;
    10'd64: brom_out <= 64'd464818087266499824;
    10'd65: brom_out <= 64'd2978682856478279174;
    10'd66: brom_out <= 64'd7468303068922238782;
    10'd67: brom_out <= 64'd4588180871198807947;
    10'd68: brom_out <= 64'd7558443736800330221;
    10'd69: brom_out <= 64'd7858840650730206709;
    10'd70: brom_out <= 64'd3151325858749743622;
    10'd71: brom_out <= 64'd3928240924200250960;
    10'd72: brom_out <= 64'd8736971688408295688;
    10'd73: brom_out <= 64'd2963845791636337106;
    10'd74: brom_out <= 64'd8638275777585364049;
    10'd75: brom_out <= 64'd4424908658087577485;
    10'd76: brom_out <= 64'd3711910516821046543;
    10'd77: brom_out <= 64'd564452646185648433;
    10'd78: brom_out <= 64'd351604139475031744;
    10'd79: brom_out <= 64'd3218941757365961417;
    10'd80: brom_out <= 64'd3971250007542337134;
    10'd81: brom_out <= 64'd6348148117183227029;
    10'd82: brom_out <= 64'd6375967769309133740;
    10'd83: brom_out <= 64'd2697116720289292087;
    10'd84: brom_out <= 64'd6627704934952898664;
    10'd85: brom_out <= 64'd3922405524646050047;
    10'd86: brom_out <= 64'd9046808849552815412;
    10'd87: brom_out <= 64'd8034888508511925711;
    10'd88: brom_out <= 64'd2859666381547961291;
    10'd89: brom_out <= 64'd7137160280198859230;
    10'd90: brom_out <= 64'd8110123499042701751;
    10'd91: brom_out <= 64'd8034333698633526839;
    10'd92: brom_out <= 64'd4803581755516584292;
    10'd93: brom_out <= 64'd4590259300347101331;
    10'd94: brom_out <= 64'd1559091360608078193;
    10'd95: brom_out <= 64'd1403053605871108975;
    10'd96: brom_out <= 64'd4595273378699324055;
    10'd97: brom_out <= 64'd2776148100713341227;
    10'd98: brom_out <= 64'd2594924969993574608;
    10'd99: brom_out <= 64'd7071793234846935066;
    10'd100: brom_out <= 64'd2462386169309760855;
    10'd101: brom_out <= 64'd3231532715502928322;
    10'd102: brom_out <= 64'd9198317650626931837;
    10'd103: brom_out <= 64'd4609249902052002620;
    10'd104: brom_out <= 64'd7549026117124348284;
    10'd105: brom_out <= 64'd7171373982066933827;
    10'd106: brom_out <= 64'd5368887724683895641;
    10'd107: brom_out <= 64'd4062746511325342569;
    10'd108: brom_out <= 64'd7171535623464460640;
    10'd109: brom_out <= 64'd7741372681338336922;
    10'd110: brom_out <= 64'd3162624206701104350;
    10'd111: brom_out <= 64'd855955066017895617;
    10'd112: brom_out <= 64'd1930668069630434611;
    10'd113: brom_out <= 64'd2928098416169300648;
    10'd114: brom_out <= 64'd5854960979430630462;
    10'd115: brom_out <= 64'd5811220473517558745;
    10'd116: brom_out <= 64'd1456145562961886765;
    10'd117: brom_out <= 64'd4416594423745725139;
    10'd118: brom_out <= 64'd2376547190173544320;
    10'd119: brom_out <= 64'd5727465189061744601;
    10'd120: brom_out <= 64'd7788324255361591123;
    10'd121: brom_out <= 64'd6767070414593594546;
    10'd122: brom_out <= 64'd6186496404391441263;
    10'd123: brom_out <= 64'd3140361231570247381;
    10'd124: brom_out <= 64'd8400656207709953750;
    10'd125: brom_out <= 64'd7036353943044608377;
    10'd126: brom_out <= 64'd5075091738590864952;
    10'd127: brom_out <= 64'd2397774606766741304;
    10'd128: brom_out <= 64'd6226365014916112750;
    10'd129: brom_out <= 64'd5428798789970012252;
    10'd130: brom_out <= 64'd5439353873355781496;
    10'd131: brom_out <= 64'd5571426184817407302;
    10'd132: brom_out <= 64'd1969591382671456713;
    10'd133: brom_out <= 64'd5181737157734702211;
    10'd134: brom_out <= 64'd7892990332141014012;
    10'd135: brom_out <= 64'd6159890351897691019;
    10'd136: brom_out <= 64'd1003510499900998868;
    10'd137: brom_out <= 64'd2671016986383601893;
    10'd138: brom_out <= 64'd3143394533206848762;
    10'd139: brom_out <= 64'd695344718632048640;
    10'd140: brom_out <= 64'd7053302599317773964;
    10'd141: brom_out <= 64'd1699346888481008308;
    10'd142: brom_out <= 64'd2698649976683576475;
    10'd143: brom_out <= 64'd7401947428770721099;
    10'd144: brom_out <= 64'd5933913752163124397;
    10'd145: brom_out <= 64'd5935407879197926157;
    10'd146: brom_out <= 64'd2993336536115385941;
    10'd147: brom_out <= 64'd55271682771906773;
    10'd148: brom_out <= 64'd8676893857881770324;
    10'd149: brom_out <= 64'd1518683083191258302;
    10'd150: brom_out <= 64'd8936281099231278912;
    10'd151: brom_out <= 64'd3525165000835027303;
    10'd152: brom_out <= 64'd4684591512257835936;
    10'd153: brom_out <= 64'd3370585482942522412;
    10'd154: brom_out <= 64'd5026403576168103312;
    10'd155: brom_out <= 64'd5048938432560231129;
    10'd156: brom_out <= 64'd4821552287445869606;
    10'd157: brom_out <= 64'd3812697702688826811;
    10'd158: brom_out <= 64'd849666076645434347;
    10'd159: brom_out <= 64'd7935697742826921448;
    10'd160: brom_out <= 64'd1365445091898096717;
    10'd161: brom_out <= 64'd590904085002712108;
    10'd162: brom_out <= 64'd254296121785148329;
    10'd163: brom_out <= 64'd5346302256075872931;
    10'd164: brom_out <= 64'd4054681239756612468;
    10'd165: brom_out <= 64'd983295328193775601;
    10'd166: brom_out <= 64'd3708187878323388551;
    10'd167: brom_out <= 64'd1439765824625554834;
    10'd168: brom_out <= 64'd171317774340299743;
    10'd169: brom_out <= 64'd3342451613070614823;
    10'd170: brom_out <= 64'd5541098046248861058;
    10'd171: brom_out <= 64'd1186113301195529614;
    10'd172: brom_out <= 64'd315448615540709982;
    10'd173: brom_out <= 64'd6365930435172523419;
    10'd174: brom_out <= 64'd4153742913801987991;
    10'd175: brom_out <= 64'd2331867165497853675;
    10'd176: brom_out <= 64'd6872169185807671677;
    10'd177: brom_out <= 64'd1232811821993946514;
    10'd178: brom_out <= 64'd1246495513601107867;
    10'd179: brom_out <= 64'd3765133689885438821;
    10'd180: brom_out <= 64'd6217630793046153812;
    10'd181: brom_out <= 64'd2957561813401634546;
    10'd182: brom_out <= 64'd4181500022422225997;
    10'd183: brom_out <= 64'd186757822164256883;
    10'd184: brom_out <= 64'd4252343237914006313;
    10'd185: brom_out <= 64'd2167868220626469006;
    10'd186: brom_out <= 64'd642809596208760966;
    10'd187: brom_out <= 64'd5132149445250676656;
    10'd188: brom_out <= 64'd5047811918853047176;
    10'd189: brom_out <= 64'd3681996519355107202;
    10'd190: brom_out <= 64'd2062831261923496231;
    10'd191: brom_out <= 64'd2070164934788009753;
    10'd192: brom_out <= 64'd7089614964709898385;
    10'd193: brom_out <= 64'd99797742496628440;
    10'd194: brom_out <= 64'd93597724244979478;
    10'd195: brom_out <= 64'd2703188527959273500;
    10'd196: brom_out <= 64'd525111339311974560;
    10'd197: brom_out <= 64'd2073887859079328870;
    10'd198: brom_out <= 64'd7010507675909334974;
    10'd199: brom_out <= 64'd5071654422350367605;
    10'd200: brom_out <= 64'd542861560934892170;
    10'd201: brom_out <= 64'd8260504402447994528;
    10'd202: brom_out <= 64'd6292353272454494027;
    10'd203: brom_out <= 64'd4470779827374382672;
    10'd204: brom_out <= 64'd2903936630100625707;
    10'd205: brom_out <= 64'd457501523175826886;
    10'd206: brom_out <= 64'd3954015878074795233;
    10'd207: brom_out <= 64'd8008368157905688049;
    10'd208: brom_out <= 64'd1057877703198774963;
    10'd209: brom_out <= 64'd7321797862192810070;
    10'd210: brom_out <= 64'd881446925189189622;
    10'd211: brom_out <= 64'd6180881228235604727;
    10'd212: brom_out <= 64'd5145557019096535373;
    10'd213: brom_out <= 64'd5399562539430498850;
    10'd214: brom_out <= 64'd2097536514174451427;
    10'd215: brom_out <= 64'd1302969704392912586;
    10'd216: brom_out <= 64'd6383088688177896759;
    10'd217: brom_out <= 64'd4776820405731634442;
    10'd218: brom_out <= 64'd7485706981003727294;
    10'd219: brom_out <= 64'd7218866889904024957;
    10'd220: brom_out <= 64'd5642552092961002333;
    10'd221: brom_out <= 64'd6355105950674987139;
    10'd222: brom_out <= 64'd7444903694469134013;
    10'd223: brom_out <= 64'd6656058382601779780;
    10'd224: brom_out <= 64'd5716724314729095879;
    10'd225: brom_out <= 64'd7516010632001644383;
    10'd226: brom_out <= 64'd1761043349758399802;
    10'd227: brom_out <= 64'd8728872155849937065;
    10'd228: brom_out <= 64'd3572156180491922781;
    10'd229: brom_out <= 64'd1535975523511082697;
    10'd230: brom_out <= 64'd2643693107760143504;
    10'd231: brom_out <= 64'd6280050499334699438;
    10'd232: brom_out <= 64'd3478111344349331952;
    10'd233: brom_out <= 64'd9205850204399306455;
    10'd234: brom_out <= 64'd1782213838681283426;
    10'd235: brom_out <= 64'd828337951715771591;
    10'd236: brom_out <= 64'd6445385301812469258;
    10'd237: brom_out <= 64'd1475549944326657173;
    10'd238: brom_out <= 64'd4471481750525228472;
    10'd239: brom_out <= 64'd7756338194758556395;
    10'd240: brom_out <= 64'd8889570641836897678;
    10'd241: brom_out <= 64'd9214805754961653984;
    10'd242: brom_out <= 64'd7744392375168708057;
    10'd243: brom_out <= 64'd2777060205167971659;
    10'd244: brom_out <= 64'd4498277668647537036;
    10'd245: brom_out <= 64'd218799722747709959;
    10'd246: brom_out <= 64'd6191163825205153709;
    10'd247: brom_out <= 64'd2748131089998747006;
    10'd248: brom_out <= 64'd7096711168948612233;
    10'd249: brom_out <= 64'd1406004993547085630;
    10'd250: brom_out <= 64'd6104292625726894888;
    10'd251: brom_out <= 64'd4919191232943017838;
    10'd252: brom_out <= 64'd5368845909558099263;
    10'd253: brom_out <= 64'd295428738034846021;
    10'd254: brom_out <= 64'd2308711598608464189;
    10'd255: brom_out <= 64'd6096319519375431872;
    10'd256: brom_out <= 64'd6192068958546582061;
    10'd257: brom_out <= 64'd1159693055014920082;
    10'd258: brom_out <= 64'd1796322016343730656;
    10'd259: brom_out <= 64'd125741342203844633;
    10'd260: brom_out <= 64'd7272549208785566368;
    10'd261: brom_out <= 64'd3305972630871509593;
    10'd262: brom_out <= 64'd7788251043344017392;
    10'd263: brom_out <= 64'd7754941374064063869;
    10'd264: brom_out <= 64'd7150486235490755525;
    10'd265: brom_out <= 64'd5572229739443640910;
    10'd266: brom_out <= 64'd7237377075799460817;
    10'd267: brom_out <= 64'd7262655534050751425;
    10'd268: brom_out <= 64'd2039786129721060611;
    10'd269: brom_out <= 64'd2897246424902218592;
    10'd270: brom_out <= 64'd2721707540031427017;
    10'd271: brom_out <= 64'd5113335136394915301;
    10'd272: brom_out <= 64'd6726333986398514634;
    10'd273: brom_out <= 64'd5879912706154820525;
    10'd274: brom_out <= 64'd710295836467163914;
    10'd275: brom_out <= 64'd5469361348601251500;
    10'd276: brom_out <= 64'd7220067846396189031;
    10'd277: brom_out <= 64'd7533447111696801148;
    10'd278: brom_out <= 64'd2145807780165639437;
    10'd279: brom_out <= 64'd9105128469287532002;
    10'd280: brom_out <= 64'd3514511250914930670;
    10'd281: brom_out <= 64'd7719981404049964815;
    10'd282: brom_out <= 64'd4609468238257219661;
    10'd283: brom_out <= 64'd1693288256086857860;
    10'd284: brom_out <= 64'd1937057571872129234;
    10'd285: brom_out <= 64'd1118118188210935647;
    10'd286: brom_out <= 64'd8123032552857054094;
    10'd287: brom_out <= 64'd4933353624348031646;
    10'd288: brom_out <= 64'd8509966626912802274;
    10'd289: brom_out <= 64'd5286704066961376178;
    10'd290: brom_out <= 64'd529000162962455889;
    10'd291: brom_out <= 64'd1060530080179134359;
    10'd292: brom_out <= 64'd7885391976349690460;
    10'd293: brom_out <= 64'd4704030701995566024;
    10'd294: brom_out <= 64'd5941448696335591560;
    10'd295: brom_out <= 64'd8343321056375228956;
    10'd296: brom_out <= 64'd5740388156642824243;
    10'd297: brom_out <= 64'd2741573671984257673;
    10'd298: brom_out <= 64'd4825669769055971489;
    10'd299: brom_out <= 64'd6204443521919095712;
    10'd300: brom_out <= 64'd3453819474470703498;
    10'd301: brom_out <= 64'd6519975654949489323;
    10'd302: brom_out <= 64'd3465890630705710859;
    10'd303: brom_out <= 64'd1636504433951697239;
    10'd304: brom_out <= 64'd3160378248132958205;
    10'd305: brom_out <= 64'd8079195116669884562;
    10'd306: brom_out <= 64'd1330718716890237459;
    10'd307: brom_out <= 64'd5981615816055793875;
    10'd308: brom_out <= 64'd8498120993252165605;
    10'd309: brom_out <= 64'd7710571130249687669;
    10'd310: brom_out <= 64'd8433949220284074317;
    10'd311: brom_out <= 64'd7891691529848080392;
    10'd312: brom_out <= 64'd6814828678859471793;
    10'd313: brom_out <= 64'd4007664876865617149;
    10'd314: brom_out <= 64'd3904923598349859840;
    10'd315: brom_out <= 64'd6360480171627733212;
    10'd316: brom_out <= 64'd2309708901247373513;
    10'd317: brom_out <= 64'd1525121092500310936;
    10'd318: brom_out <= 64'd16669355320858615;
    10'd319: brom_out <= 64'd5930297400455869884;
    10'd320: brom_out <= 64'd8393046322456432693;
    10'd321: brom_out <= 64'd5590106815304323809;
    10'd322: brom_out <= 64'd782535549554235096;
    10'd323: brom_out <= 64'd2633259836156076026;
    10'd324: brom_out <= 64'd5777401271193676712;
    10'd325: brom_out <= 64'd9027064800603781502;
    10'd326: brom_out <= 64'd8550452487403366270;
    10'd327: brom_out <= 64'd5166206035685481241;
    10'd328: brom_out <= 64'd7808713511810165244;
    10'd329: brom_out <= 64'd274459991172651778;
    10'd330: brom_out <= 64'd910815956873772067;
    10'd331: brom_out <= 64'd3037646691043026641;
    10'd332: brom_out <= 64'd4545698443082775269;
    10'd333: brom_out <= 64'd2454827340098860676;
    10'd334: brom_out <= 64'd3511687562711658340;
    10'd335: brom_out <= 64'd5372332410628907647;
    10'd336: brom_out <= 64'd2903391995836245846;
    10'd337: brom_out <= 64'd7231088699097087118;
    10'd338: brom_out <= 64'd549751111443322344;
    10'd339: brom_out <= 64'd2285120989557309564;
    10'd340: brom_out <= 64'd8403344402217028520;
    10'd341: brom_out <= 64'd7807489848643099872;
    10'd342: brom_out <= 64'd3230936237772476709;
    10'd343: brom_out <= 64'd1826597817821362425;
    10'd344: brom_out <= 64'd1772554492871977253;
    10'd345: brom_out <= 64'd2703486256765177688;
    10'd346: brom_out <= 64'd6074570912297676648;
    10'd347: brom_out <= 64'd8527702417501121898;
    10'd348: brom_out <= 64'd4439316959389010555;
    10'd349: brom_out <= 64'd4457589562422976492;
    10'd350: brom_out <= 64'd1686195917870897324;
    10'd351: brom_out <= 64'd2634402486982227113;
    10'd352: brom_out <= 64'd8311611936398516071;
    10'd353: brom_out <= 64'd4589438600012943360;
    10'd354: brom_out <= 64'd2939837104655752758;
    10'd355: brom_out <= 64'd4114796635571823452;
    10'd356: brom_out <= 64'd5464798183059646670;
    10'd357: brom_out <= 64'd1088054060805478255;
    10'd358: brom_out <= 64'd791846980082136773;
    10'd359: brom_out <= 64'd3475654310643013931;
    10'd360: brom_out <= 64'd474952354993185951;
    10'd361: brom_out <= 64'd5006024000541207715;
    10'd362: brom_out <= 64'd384653518295825934;
    10'd363: brom_out <= 64'd4102273044726344936;
    10'd364: brom_out <= 64'd5092186480685169789;
    10'd365: brom_out <= 64'd970407159055326691;
    10'd366: brom_out <= 64'd8416600520250423393;
    10'd367: brom_out <= 64'd3811956848453683394;
    10'd368: brom_out <= 64'd3802174757001909501;
    10'd369: brom_out <= 64'd5716198678405800318;
    10'd370: brom_out <= 64'd6613004936743467885;
    10'd371: brom_out <= 64'd6704070386751638137;
    10'd372: brom_out <= 64'd9131384685250673047;
    10'd373: brom_out <= 64'd6418341525623774333;
    10'd374: brom_out <= 64'd6083936184710043655;
    10'd375: brom_out <= 64'd3653762495492708470;
    10'd376: brom_out <= 64'd671734621348727751;
    10'd377: brom_out <= 64'd7683742792227989990;
    10'd378: brom_out <= 64'd3658421000540823124;
    10'd379: brom_out <= 64'd4374531459368300331;
    10'd380: brom_out <= 64'd3481243893374645815;
    10'd381: brom_out <= 64'd6423834149750828846;
    10'd382: brom_out <= 64'd6496458060619864987;
    10'd383: brom_out <= 64'd73115702428814728;
    10'd384: brom_out <= 64'd5092893496853917981;
    10'd385: brom_out <= 64'd8104779419146586040;
    10'd386: brom_out <= 64'd2629450283998933562;
    10'd387: brom_out <= 64'd3447848646533986482;
    10'd388: brom_out <= 64'd3041491119357596756;
    10'd389: brom_out <= 64'd5590006942133622896;
    10'd390: brom_out <= 64'd3677685952189080387;
    10'd391: brom_out <= 64'd5356739564702495632;
    10'd392: brom_out <= 64'd851648653200964577;
    10'd393: brom_out <= 64'd3062872915943182163;
    10'd394: brom_out <= 64'd4900660886885495029;
    10'd395: brom_out <= 64'd5898954515569430162;
    10'd396: brom_out <= 64'd7615771091702393585;
    10'd397: brom_out <= 64'd4672078910986180009;
    10'd398: brom_out <= 64'd1770852207371354959;
    10'd399: brom_out <= 64'd5004739783656384059;
    10'd400: brom_out <= 64'd7183136206197164704;
    10'd401: brom_out <= 64'd2082649850366603233;
    10'd402: brom_out <= 64'd5754960465788828671;
    10'd403: brom_out <= 64'd8126030331689327503;
    10'd404: brom_out <= 64'd3674101832191375914;
    10'd405: brom_out <= 64'd8436031112007516294;
    10'd406: brom_out <= 64'd3420724527339245397;
    10'd407: brom_out <= 64'd2971042736389827617;
    10'd408: brom_out <= 64'd5354840259809471406;
    10'd409: brom_out <= 64'd6502030931363910012;
    10'd410: brom_out <= 64'd8082335182850891239;
    10'd411: brom_out <= 64'd6891379871979469209;
    10'd412: brom_out <= 64'd405907765057076070;
    10'd413: brom_out <= 64'd887049970650210440;
    10'd414: brom_out <= 64'd3816324442758772072;
    10'd415: brom_out <= 64'd6289362640447157950;
    10'd416: brom_out <= 64'd6418908070461903066;
    10'd417: brom_out <= 64'd5749584372316613521;
    10'd418: brom_out <= 64'd2921731644866569442;
    10'd419: brom_out <= 64'd1238162031325735639;
    10'd420: brom_out <= 64'd6112153388438338429;
    10'd421: brom_out <= 64'd8009637371351193764;
    10'd422: brom_out <= 64'd8244651509728621613;
    10'd423: brom_out <= 64'd1106004145925981652;
    10'd424: brom_out <= 64'd7850002919444789231;
    10'd425: brom_out <= 64'd2427144979182931677;
    10'd426: brom_out <= 64'd905783496647377649;
    10'd427: brom_out <= 64'd5707305389422039546;
    10'd428: brom_out <= 64'd627693652887958811;
    10'd429: brom_out <= 64'd2086194074522431943;
    10'd430: brom_out <= 64'd6059762108987520627;
    10'd431: brom_out <= 64'd7814684497170443018;
    10'd432: brom_out <= 64'd8932176433010955680;
    10'd433: brom_out <= 64'd6375058431913780216;
    10'd434: brom_out <= 64'd5169358040688764590;
    10'd435: brom_out <= 64'd8358103728168199685;
    10'd436: brom_out <= 64'd4324478860236046205;
    10'd437: brom_out <= 64'd2297341559366227789;
    10'd438: brom_out <= 64'd2612561540033688125;
    10'd439: brom_out <= 64'd876497314882415696;
    10'd440: brom_out <= 64'd2196127990188231199;
    10'd441: brom_out <= 64'd227630122870199807;
    10'd442: brom_out <= 64'd4428649042435799499;
    10'd443: brom_out <= 64'd2916704459885367771;
    10'd444: brom_out <= 64'd5893549336767137602;
    10'd445: brom_out <= 64'd700378874414762158;
    10'd446: brom_out <= 64'd4711006633192894016;
    10'd447: brom_out <= 64'd6658948292127782393;
    10'd448: brom_out <= 64'd8577074918757021325;
    10'd449: brom_out <= 64'd5566332270607767372;
    10'd450: brom_out <= 64'd1245261505811658328;
    10'd451: brom_out <= 64'd4437855641101196385;
    10'd452: brom_out <= 64'd5403327744443637485;
    10'd453: brom_out <= 64'd1998936166749516770;
    10'd454: brom_out <= 64'd4637437027325163928;
    10'd455: brom_out <= 64'd1820109539653306332;
    10'd456: brom_out <= 64'd1238821654401532501;
    10'd457: brom_out <= 64'd9012166713295197499;
    10'd458: brom_out <= 64'd4140196495551771412;
    10'd459: brom_out <= 64'd4708243363225416979;
    10'd460: brom_out <= 64'd7678697812724703979;
    10'd461: brom_out <= 64'd1942794318847553323;
    10'd462: brom_out <= 64'd7513766008916832273;
    10'd463: brom_out <= 64'd3956455137604811437;
    10'd464: brom_out <= 64'd3474109625556721727;
    10'd465: brom_out <= 64'd9175631247054802132;
    10'd466: brom_out <= 64'd8587516205661733991;
    10'd467: brom_out <= 64'd2730435499985491472;
    10'd468: brom_out <= 64'd8266806500775076411;
    10'd469: brom_out <= 64'd2765582965792247542;
    10'd470: brom_out <= 64'd87548571312450736;
    10'd471: brom_out <= 64'd6338855802636615286;
    10'd472: brom_out <= 64'd4331841088716863106;
    10'd473: brom_out <= 64'd7370417326155807593;
    10'd474: brom_out <= 64'd2708856365737743494;
    10'd475: brom_out <= 64'd522163652426224221;
    10'd476: brom_out <= 64'd3957354033542795518;
    10'd477: brom_out <= 64'd4070727811731289008;
    10'd478: brom_out <= 64'd7777763553641271790;
    10'd479: brom_out <= 64'd6949754382192805521;
    10'd480: brom_out <= 64'd6284107821877667060;
    10'd481: brom_out <= 64'd597411352177070931;
    10'd482: brom_out <= 64'd6164721133495571031;
    10'd483: brom_out <= 64'd5570579181901818869;
    10'd484: brom_out <= 64'd2941157606459076432;
    10'd485: brom_out <= 64'd2175496214153705066;
    10'd486: brom_out <= 64'd6086604863266952663;
    10'd487: brom_out <= 64'd4708479177706903053;
    10'd488: brom_out <= 64'd5408360093042724747;
    10'd489: brom_out <= 64'd2583084939302978673;
    10'd490: brom_out <= 64'd3827754383887830875;
    10'd491: brom_out <= 64'd6987828419030564022;
    10'd492: brom_out <= 64'd8585572637166925618;
    10'd493: brom_out <= 64'd2871615205384557091;
    10'd494: brom_out <= 64'd2279506272437617033;
    10'd495: brom_out <= 64'd2466579790451595447;
    10'd496: brom_out <= 64'd5610224495861148711;
    10'd497: brom_out <= 64'd4655293031232142642;
    10'd498: brom_out <= 64'd967077408856567116;
    10'd499: brom_out <= 64'd974279068567969527;
    10'd500: brom_out <= 64'd4535950713114274704;
    10'd501: brom_out <= 64'd8675110334873814678;
    10'd502: brom_out <= 64'd119908315201321689;
    10'd503: brom_out <= 64'd724891155700559232;
    10'd504: brom_out <= 64'd1333660446184381421;
    10'd505: brom_out <= 64'd7833308126742092808;
    10'd506: brom_out <= 64'd2796274755128593469;
    10'd507: brom_out <= 64'd77184575555698474;
    10'd508: brom_out <= 64'd2091401977497967068;
    10'd509: brom_out <= 64'd2479352029885404790;
    10'd510: brom_out <= 64'd934841504910444507;
    10'd511: brom_out <= 64'd3210500733866020013;
    default: brom_out <= 64'h1;
    endcase
end

generate
    if(DELAY == 1) begin
        assign b = brom_out;
    end
endgenerate

endmodule

//-------------------------------------------------------------------------------------------------

module tw_rom_10_intt_nwc
#(
    parameter LOGN  = 10,
    parameter LOGQ  = 64,
    parameter DELAY = 1,
    parameter STAGE = 10
)(
    input            clk,
    input [LOGN-1:0] raddr,
    output[LOGQ-1:0] b
);

(* ram_style = "block" *)
reg [LOGQ-1:0] brom_out, brom_out2;

always @(posedge clk) begin
    case(raddr[STAGE-1:0])
    11'd0: brom_out <= 64'd155299545700672449;
    11'd1: brom_out <= 64'd8591586975124194640;
    11'd2: brom_out <= 64'd3167401383237838777;
    11'd3: brom_out <= 64'd591188586763527378;
    11'd4: brom_out <= 64'd1514599663756940472;
    11'd5: brom_out <= 64'd7817930662417897360;
    11'd6: brom_out <= 64'd3620991004643695475;
    11'd7: brom_out <= 64'd7542692879326719854;
    11'd8: brom_out <= 64'd7902824838328275304;
    11'd9: brom_out <= 64'd763189247563564006;
    11'd10: brom_out <= 64'd8774968117827411067;
    11'd11: brom_out <= 64'd7673518914872814072;
    11'd12: brom_out <= 64'd5373092361287203993;
    11'd13: brom_out <= 64'd3876460951776019299;
    11'd14: brom_out <= 64'd4760195863663172767;
    11'd15: brom_out <= 64'd548897859864734688;
    11'd16: brom_out <= 64'd8908024222468824634;
    11'd17: brom_out <= 64'd5928464271996740273;
    11'd18: brom_out <= 64'd5908873892802598358;
    11'd19: brom_out <= 64'd1780406181529146949;
    11'd20: brom_out <= 64'd5736893487197545155;
    11'd21: brom_out <= 64'd2356070081099186446;
    11'd22: brom_out <= 64'd1418818644174705489;
    11'd23: brom_out <= 64'd2084377973795870866;
    11'd24: brom_out <= 64'd6144362497601089118;
    11'd25: brom_out <= 64'd7123992511842491259;
    11'd26: brom_out <= 64'd4466959297753725853;
    11'd27: brom_out <= 64'd915255655171031995;
    11'd28: brom_out <= 64'd412784429296323548;
    11'd29: brom_out <= 64'd2607976344674075427;
    11'd30: brom_out <= 64'd3806348048038220265;
    11'd31: brom_out <= 64'd3627078416448126394;
    11'd32: brom_out <= 64'd1158029312224390638;
    11'd33: brom_out <= 64'd8529432223335041238;
    11'd34: brom_out <= 64'd6055478084367806153;
    11'd35: brom_out <= 64'd1522346900703918240;
    11'd36: brom_out <= 64'd2943964933625184572;
    11'd37: brom_out <= 64'd6279056307255967124;
    11'd38: brom_out <= 64'd1310717603008154032;
    11'd39: brom_out <= 64'd2036871276625425044;
    11'd40: brom_out <= 64'd549090306655750826;
    11'd41: brom_out <= 64'd8254812355918294849;
    11'd42: brom_out <= 64'd3751939551327780519;
    11'd43: brom_out <= 64'd4700199910743006656;
    11'd44: brom_out <= 64'd7651159289997704313;
    11'd45: brom_out <= 64'd6174118643639414798;
    11'd46: brom_out <= 64'd1821201232213099039;
    11'd47: brom_out <= 64'd7549080415689794490;
    11'd48: brom_out <= 64'd4134920192217805033;
    11'd49: brom_out <= 64'd1566244339874456380;
    11'd50: brom_out <= 64'd8941755252885023556;
    11'd51: brom_out <= 64'd8259111416425220548;
    11'd52: brom_out <= 64'd6863892824799961069;
    11'd53: brom_out <= 64'd4094211991695582914;
    11'd54: brom_out <= 64'd1017338174540963918;
    11'd55: brom_out <= 64'd8231638915758483851;
    11'd56: brom_out <= 64'd1545147831700695205;
    11'd57: brom_out <= 64'd6286107393354575151;
    11'd58: brom_out <= 64'd866731065849342802;
    11'd59: brom_out <= 64'd5817704039855958750;
    11'd60: brom_out <= 64'd1144960696522762897;
    11'd61: brom_out <= 64'd3079619532358567389;
    11'd62: brom_out <= 64'd3641446469606875086;
    11'd63: brom_out <= 64'd4849465172743338905;
    11'd64: brom_out <= 64'd9198110032305492864;
    11'd65: brom_out <= 64'd8935961102750503989;
    11'd66: brom_out <= 64'd7338214287406543596;
    11'd67: brom_out <= 64'd6144254994690576277;
    11'd68: brom_out <= 64'd8070099755377702019;
    11'd69: brom_out <= 64'd4610586010050803807;
    11'd70: brom_out <= 64'd6317856931341908110;
    11'd71: brom_out <= 64'd1836558788137277687;
    11'd72: brom_out <= 64'd5391618511616287733;
    11'd73: brom_out <= 64'd7807583818559962560;
    11'd74: brom_out <= 64'd3178626018632929050;
    11'd75: brom_out <= 64'd6077672357582230492;
    11'd76: brom_out <= 64'd1609504591888863414;
    11'd77: brom_out <= 64'd1103508469039991957;
    11'd78: brom_out <= 64'd1642907077317613831;
    11'd79: brom_out <= 64'd4007859166999782559;
    11'd80: brom_out <= 64'd7508353885558613582;
    11'd81: brom_out <= 64'd4364643021443062444;
    11'd82: brom_out <= 64'd7703804984359951860;
    11'd83: brom_out <= 64'd5273994222492752369;
    11'd84: brom_out <= 64'd5578329071142226718;
    11'd85: brom_out <= 64'd7430686175918402487;
    11'd86: brom_out <= 64'd2509304031536307347;
    11'd87: brom_out <= 64'd477446785469947360;
    11'd88: brom_out <= 64'd6477068066809356990;
    11'd89: brom_out <= 64'd8031446026159174764;
    11'd90: brom_out <= 64'd2687264344494152543;
    11'd91: brom_out <= 64'd6581341717046937685;
    11'd92: brom_out <= 64'd4639658250367395091;
    11'd93: brom_out <= 64'd3891637693217679590;
    11'd94: brom_out <= 64'd1059820646701210258;
    11'd95: brom_out <= 64'd818722698256349410;
    11'd96: brom_out <= 64'd4049312626161446516;
    11'd97: brom_out <= 64'd3004162438510806775;
    11'd98: brom_out <= 64'd6784195684454936881;
    11'd99: brom_out <= 64'd5404780470263141518;
    11'd100: brom_out <= 64'd819871369487893246;
    11'd101: brom_out <= 64'd6183641390300895460;
    11'd102: brom_out <= 64'd8614975202109589732;
    11'd103: brom_out <= 64'd4968747041835250263;
    11'd104: brom_out <= 64'd7323236899119000345;
    11'd105: brom_out <= 64'd6327047866211201412;
    11'd106: brom_out <= 64'd6303414007022090464;
    11'd107: brom_out <= 64'd7566815562484798677;
    11'd108: brom_out <= 64'd6901929863486149509;
    11'd109: brom_out <= 64'd8222690866176161287;
    11'd110: brom_out <= 64'd2522460457842332837;
    11'd111: brom_out <= 64'd4220581074784152971;
    11'd112: brom_out <= 64'd6238879527834839958;
    11'd113: brom_out <= 64'd919631675990915272;
    11'd114: brom_out <= 64'd5519785635586850819;
    11'd115: brom_out <= 64'd8208831059893882519;
    11'd116: brom_out <= 64'd4915421594627397633;
    11'd117: brom_out <= 64'd7586062489076878287;
    11'd118: brom_out <= 64'd7617204530614757254;
    11'd119: brom_out <= 64'd1070383556442660744;
    11'd120: brom_out <= 64'd8140858962325166315;
    11'd121: brom_out <= 64'd4908397430704463857;
    11'd122: brom_out <= 64'd6980561833182397069;
    11'd123: brom_out <= 64'd8028669790929027125;
    11'd124: brom_out <= 64'd8580458598856579249;
    11'd125: brom_out <= 64'd3216346525908124941;
    11'd126: brom_out <= 64'd3832635110383635309;
    11'd127: brom_out <= 64'd5274665080719022868;
    11'd128: brom_out <= 64'd761644425330199272;
    11'd129: brom_out <= 64'd2991460051583178365;
    11'd130: brom_out <= 64'd706928156095515790;
    11'd131: brom_out <= 64'd8254874734866087170;
    11'd132: brom_out <= 64'd4579564535757996383;
    11'd133: brom_out <= 64'd4994771842306729102;
    11'd134: brom_out <= 64'd9187349396686375108;
    11'd135: brom_out <= 64'd1250536128227672786;
    11'd136: brom_out <= 64'd2519346554143507611;
    11'd137: brom_out <= 64'd5359207005777685074;
    11'd138: brom_out <= 64'd6772576518519916947;
    11'd139: brom_out <= 64'd495084928218723803;
    11'd140: brom_out <= 64'd8626187869693540491;
    11'd141: brom_out <= 64'd7636919348751616120;
    11'd142: brom_out <= 64'd3023092419124062753;
    11'd143: brom_out <= 64'd4872935445130040668;
    11'd144: brom_out <= 64'd5485806031066447759;
    11'd145: brom_out <= 64'd5407652607953428448;
    11'd146: brom_out <= 64'd4382121046488924351;
    11'd147: brom_out <= 64'd7637944378401354825;
    11'd148: brom_out <= 64'd3636639398006559632;
    11'd149: brom_out <= 64'd6230337823244594242;
    11'd150: brom_out <= 64'd1945442526511340058;
    11'd151: brom_out <= 64'd6372242758954669061;
    11'd152: brom_out <= 64'd4124955256152859363;
    11'd153: brom_out <= 64'd3126938990396619728;
    11'd154: brom_out <= 64'd1515533781493865721;
    11'd155: brom_out <= 64'd5114376596938491811;
    11'd156: brom_out <= 64'd4019065279918376385;
    11'd157: brom_out <= 64'd2369822980812815061;
    11'd158: brom_out <= 64'd4127230542017488573;
    11'd159: brom_out <= 64'd8679545142051594119;
    11'd160: brom_out <= 64'd1960525529548210299;
    11'd161: brom_out <= 64'd6068989862395001591;
    11'd162: brom_out <= 64'd6085765700274220889;
    11'd163: brom_out <= 64'd3401668953812010006;
    11'd164: brom_out <= 64'd7637335644243982898;
    11'd165: brom_out <= 64'd7483539404139064850;
    11'd166: brom_out <= 64'd1211022569296579482;
    11'd167: brom_out <= 64'd5632876105105940994;
    11'd168: brom_out <= 64'd6103576109977111487;
    11'd169: brom_out <= 64'd2318854527119863408;
    11'd170: brom_out <= 64'd1695176741447732168;
    11'd171: brom_out <= 64'd1790195042493211624;
    11'd172: brom_out <= 64'd2842565075093397561;
    11'd173: brom_out <= 64'd5435963472951530096;
    11'd174: brom_out <= 64'd5208588277951337540;
    11'd175: brom_out <= 64'd4236251210736797742;
    11'd176: brom_out <= 64'd843199340190868878;
    11'd177: brom_out <= 64'd1092512432296708951;
    11'd178: brom_out <= 64'd2946132479941139089;
    11'd179: brom_out <= 64'd7670897235897672237;
    11'd180: brom_out <= 64'd3637138387601219284;
    11'd181: brom_out <= 64'd4642477032133592860;
    11'd182: brom_out <= 64'd575745599961146758;
    11'd183: brom_out <= 64'd2793234862260117914;
    11'd184: brom_out <= 64'd7657659146000242080;
    11'd185: brom_out <= 64'd6372094233712387000;
    11'd186: brom_out <= 64'd6176174963711788051;
    11'd187: brom_out <= 64'd2319329316203352609;
    11'd188: brom_out <= 64'd6049587548814090897;
    11'd189: brom_out <= 64'd9007215134378364274;
    11'd190: brom_out <= 64'd3207576084825550941;
    11'd191: brom_out <= 64'd4202885042285007382;
    11'd192: brom_out <= 64'd2884224422498108059;
    11'd193: brom_out <= 64'd6183853536836250528;
    11'd194: brom_out <= 64'd2670454142491632319;
    11'd195: brom_out <= 64'd2320029118861391477;
    11'd196: brom_out <= 64'd8376561785798592285;
    11'd197: brom_out <= 64'd2992583618867802019;
    11'd198: brom_out <= 64'd5248188609469701482;
    11'd199: brom_out <= 64'd2762518159980585286;
    11'd200: brom_out <= 64'd4295342249137175680;
    11'd201: brom_out <= 64'd7932441453988948969;
    11'd202: brom_out <= 64'd2334660456303647272;
    11'd203: brom_out <= 64'd333205755352370400;
    11'd204: brom_out <= 64'd907921074387711606;
    11'd205: brom_out <= 64'd5166365826688214535;
    11'd206: brom_out <= 64'd9025095217715156325;
    11'd207: brom_out <= 64'd2846565905266866879;
    11'd208: brom_out <= 64'd1225666943611193327;
    11'd209: brom_out <= 64'd15116887055001170;
    11'd210: brom_out <= 64'd7750614262329275312;
    11'd211: brom_out <= 64'd1904884659095357883;
    11'd212: brom_out <= 64'd6576541357640508954;
    11'd213: brom_out <= 64'd594192566179244285;
    11'd214: brom_out <= 64'd196051014340678308;
    11'd215: brom_out <= 64'd6750046039111356045;
    11'd216: brom_out <= 64'd1253061220177896022;
    11'd217: brom_out <= 64'd4693232200421745805;
    11'd218: brom_out <= 64'd6804550799754867160;
    11'd219: brom_out <= 64'd2969038553162991539;
    11'd220: brom_out <= 64'd5935254196818449959;
    11'd221: brom_out <= 64'd1905036106355650949;
    11'd222: brom_out <= 64'd1118547525326689136;
    11'd223: brom_out <= 64'd133427282067141130;
    11'd224: brom_out <= 64'd8129343517429338242;
    11'd225: brom_out <= 64'd944368318123377314;
    11'd226: brom_out <= 64'd5326022513342054649;
    11'd227: brom_out <= 64'd5984489630834845160;
    11'd228: brom_out <= 64'd7384294585376217243;
    11'd229: brom_out <= 64'd2314043236292767398;
    11'd230: brom_out <= 64'd7171334747151766070;
    11'd231: brom_out <= 64'd9209694779854938873;
    11'd232: brom_out <= 64'd8426084403847311000;
    11'd233: brom_out <= 64'd7737471128275518782;
    11'd234: brom_out <= 64'd5182789654663425165;
    11'd235: brom_out <= 64'd3038860110131058391;
    11'd236: brom_out <= 64'd6701035787418191993;
    11'd237: brom_out <= 64'd1107423090841681213;
    11'd238: brom_out <= 64'd8680765855631139946;
    11'd239: brom_out <= 64'd7746857959523985121;
    11'd240: brom_out <= 64'd7145038203562988461;
    11'd241: brom_out <= 64'd6099584987210526395;
    11'd242: brom_out <= 64'd5734319089212947416;
    11'd243: brom_out <= 64'd9184317857101729769;
    11'd244: brom_out <= 64'd8952938491005290769;
    11'd245: brom_out <= 64'd9209525668573131033;
    11'd246: brom_out <= 64'd6928109774782512045;
    11'd247: brom_out <= 64'd6301102485076257059;
    11'd248: brom_out <= 64'd2155719515733443264;
    11'd249: brom_out <= 64'd6397179018084218993;
    11'd250: brom_out <= 64'd67710781327552919;
    11'd251: brom_out <= 64'd2220341238225044662;
    11'd252: brom_out <= 64'd3197005768988671911;
    11'd253: brom_out <= 64'd2363885441477553649;
    11'd254: brom_out <= 64'd4438981546541157226;
    11'd255: brom_out <= 64'd4250450348376300205;
    11'd256: brom_out <= 64'd5680384952025565122;
    11'd257: brom_out <= 64'd4235870775706994632;
    11'd258: brom_out <= 64'd6566997680978011943;
    11'd259: brom_out <= 64'd7031686766803585650;
    11'd260: brom_out <= 64'd7441602658178457958;
    11'd261: brom_out <= 64'd587280293564159230;
    11'd262: brom_out <= 64'd8228285085251450384;
    11'd263: brom_out <= 64'd227861438240141932;
    11'd264: brom_out <= 64'd1957054919284953502;
    11'd265: brom_out <= 64'd3193109024359937421;
    11'd266: brom_out <= 64'd7341285079701911949;
    11'd267: brom_out <= 64'd7926799563598326137;
    11'd268: brom_out <= 64'd7508888402962313385;
    11'd269: brom_out <= 64'd4096452394530652644;
    11'd270: brom_out <= 64'd5417979367025186582;
    11'd271: brom_out <= 64'd1117219549235793098;
    11'd272: brom_out <= 64'd305105216848129692;
    11'd273: brom_out <= 64'd6889452513698471590;
    11'd274: brom_out <= 64'd8306230887695200469;
    11'd275: brom_out <= 64'd7877839765223129415;
    11'd276: brom_out <= 64'd1695712013653589552;
    11'd277: brom_out <= 64'd7804872488052035288;
    11'd278: brom_out <= 64'd501858554414255797;
    11'd279: brom_out <= 64'd5552517519548695450;
    11'd280: brom_out <= 64'd5901118384392698396;
    11'd281: brom_out <= 64'd1707140316774872044;
    11'd282: brom_out <= 64'd8132051213077852955;
    11'd283: brom_out <= 64'd628536434315570033;
    11'd284: brom_out <= 64'd3104751652281427870;
    11'd285: brom_out <= 64'd136310184993758523;
    11'd286: brom_out <= 64'd8852283683242620539;
    11'd287: brom_out <= 64'd8265892164849889696;
    11'd288: brom_out <= 64'd6036839688305992863;
    11'd289: brom_out <= 64'd7518421125529715847;
    11'd290: brom_out <= 64'd905880610089459061;
    11'd291: brom_out <= 64'd6483554429539231021;
    11'd292: brom_out <= 64'd4483032727014130201;
    11'd293: brom_out <= 64'd8123049477243076994;
    11'd294: brom_out <= 64'd4501035746029695362;
    11'd295: brom_out <= 64'd6003935171596987782;
    11'd296: brom_out <= 64'd4277082693891194298;
    11'd297: brom_out <= 64'd6588743782503121009;
    11'd298: brom_out <= 64'd222881655867913949;
    11'd299: brom_out <= 64'd4298288972457114646;
    11'd300: brom_out <= 64'd2466060747743623120;
    11'd301: brom_out <= 64'd215098476944587455;
    11'd302: brom_out <= 64'd5808655089357367024;
    11'd303: brom_out <= 64'd4457943904707492604;
    11'd304: brom_out <= 64'd7205668174452334545;
    11'd305: brom_out <= 64'd5974154314505877312;
    11'd306: brom_out <= 64'd7638487797572445667;
    11'd307: brom_out <= 64'd3335216815067190723;
    11'd308: brom_out <= 64'd7001890260574642730;
    11'd309: brom_out <= 64'd8642295946453124916;
    11'd310: brom_out <= 64'd5560139906224123015;
    11'd311: brom_out <= 64'd555041558694353539;
    11'd312: brom_out <= 64'd4519563697595116006;
    11'd313: brom_out <= 64'd7573991306845316380;
    11'd314: brom_out <= 64'd7881473456017877080;
    11'd315: brom_out <= 64'd1006525196979076997;
    11'd316: brom_out <= 64'd4523253709269049564;
    11'd317: brom_out <= 64'd8707254594819930941;
    11'd318: brom_out <= 64'd3241377901120040405;
    11'd319: brom_out <= 64'd7984675317219139003;
    11'd320: brom_out <= 64'd3101214915203965202;
    11'd321: brom_out <= 64'd1837387984173499890;
    11'd322: brom_out <= 64'd7834233917730301377;
    11'd323: brom_out <= 64'd2015622700673248428;
    11'd324: brom_out <= 64'd5040030845747108458;
    11'd325: brom_out <= 64'd2415938772407823212;
    11'd326: brom_out <= 64'd1433722002351993030;
    11'd327: brom_out <= 64'd6539941664781820353;
    11'd328: brom_out <= 64'd4408504617008684023;
    11'd329: brom_out <= 64'd3465261818686834369;
    11'd330: brom_out <= 64'd6713653524672007028;
    11'd331: brom_out <= 64'd5437401648693809794;
    11'd332: brom_out <= 64'd3995727708789092284;
    11'd333: brom_out <= 64'd4036127472032525531;
    11'd334: brom_out <= 64'd159198575887530223;
    11'd335: brom_out <= 64'd3036641109561738488;
    11'd336: brom_out <= 64'd343865678935493240;
    11'd337: brom_out <= 64'd6439246072166143753;
    11'd338: brom_out <= 64'd4628571125618134296;
    11'd339: brom_out <= 64'd3076493632439937520;
    11'd340: brom_out <= 64'd6664682430781220753;
    11'd341: brom_out <= 64'd4153005133628369421;
    11'd342: brom_out <= 64'd2268588113780825554;
    11'd343: brom_out <= 64'd5264887122480875761;
    11'd344: brom_out <= 64'd7372086793767004444;
    11'd345: brom_out <= 64'd5708030460374230455;
    11'd346: brom_out <= 64'd4888307838890640558;
    11'd347: brom_out <= 64'd1715234094373408718;
    11'd348: brom_out <= 64'd3211132947674934496;
    11'd349: brom_out <= 64'd2296546007350538988;
    11'd350: brom_out <= 64'd5961886057234243599;
    11'd351: brom_out <= 64'd3238725242104465219;
    11'd352: brom_out <= 64'd4546924693874029555;
    11'd353: brom_out <= 64'd8635673233040957017;
    11'd354: brom_out <= 64'd1059541674008919025;
    11'd355: brom_out <= 64'd9079413709458579446;
    11'd356: brom_out <= 64'd9100865486099282684;
    11'd357: brom_out <= 64'd6470054339417098118;
    11'd358: brom_out <= 64'd3861234640121808167;
    11'd359: brom_out <= 64'd2041897164323761649;
    11'd360: brom_out <= 64'd6282528973883425849;
    11'd361: brom_out <= 64'd4147553875257660020;
    11'd362: brom_out <= 64'd4021868810369844860;
    11'd363: brom_out <= 64'd3026190624024450633;
    11'd364: brom_out <= 64'd4040859673712721438;
    11'd365: brom_out <= 64'd5580391360694311681;
    11'd366: brom_out <= 64'd9003205404615842122;
    11'd367: brom_out <= 64'd7465868618294216802;
    11'd368: brom_out <= 64'd5925209008378466528;
    11'd369: brom_out <= 64'd2426236768536324104;
    11'd370: brom_out <= 64'd345048554160488161;
    11'd371: brom_out <= 64'd9161542714037021833;
    11'd372: brom_out <= 64'd2056881296447787458;
    11'd373: brom_out <= 64'd8637958705318879755;
    11'd374: brom_out <= 64'd5765715887113937839;
    11'd375: brom_out <= 64'd3877542420674141204;
    11'd376: brom_out <= 64'd8721937415238049120;
    11'd377: brom_out <= 64'd8891863127268636704;
    11'd378: brom_out <= 64'd2006834673636403812;
    11'd379: brom_out <= 64'd4854770072034814620;
    11'd380: brom_out <= 64'd5215912574857899194;
    11'd381: brom_out <= 64'd3083500310684001625;
    11'd382: brom_out <= 64'd1679514009156781569;
    11'd383: brom_out <= 64'd1516722928509298446;
    11'd384: brom_out <= 64'd9110296472090570993;
    11'd385: brom_out <= 64'd3569534188498493379;
    11'd386: brom_out <= 64'd2151823758199163249;
    11'd387: brom_out <= 64'd2136808689945239668;
    11'd388: brom_out <= 64'd7295909789787026847;
    11'd389: brom_out <= 64'd2920063548427700524;
    11'd390: brom_out <= 64'd7880148991479206809;
    11'd391: brom_out <= 64'd7118701410115154909;
    11'd392: brom_out <= 64'd1605173767746043079;
    11'd393: brom_out <= 64'd7055372734456367617;
    11'd394: brom_out <= 64'd1082497889398447644;
    11'd395: brom_out <= 64'd5961558258280817543;
    11'd396: brom_out <= 64'd2143166744357043707;
    11'd397: brom_out <= 64'd867574279916578313;
    11'd398: brom_out <= 64'd4410489590481103875;
    11'd399: brom_out <= 64'd4896676853699393541;
    11'd400: brom_out <= 64'd743152652173849656;
    11'd401: brom_out <= 64'd8766665715469405584;
    11'd402: brom_out <= 64'd8754802373594006508;
    11'd403: brom_out <= 64'd5163749268343386351;
    11'd404: brom_out <= 64'd808796630149307137;
    11'd405: brom_out <= 64'd5678851920497765269;
    11'd406: brom_out <= 64'd5581109811018878381;
    11'd407: brom_out <= 64'd4598202136672007123;
    11'd408: brom_out <= 64'd6717021764930164836;
    11'd409: brom_out <= 64'd3775919494807408981;
    11'd410: brom_out <= 64'd4334001442495861140;
    11'd411: brom_out <= 64'd5727022885375199616;
    11'd412: brom_out <= 64'd8607537486166103419;
    11'd413: brom_out <= 64'd2727899720984247443;
    11'd414: brom_out <= 64'd7100543299987926329;
    11'd415: brom_out <= 64'd2607449038816057334;
    11'd416: brom_out <= 64'd4106809335773449212;
    11'd417: brom_out <= 64'd5782471955832207765;
    11'd418: brom_out <= 64'd1023817687677161595;
    11'd419: brom_out <= 64'd1701747638390805703;
    11'd420: brom_out <= 64'd6701950431810787774;
    11'd421: brom_out <= 64'd8358951084842755944;
    11'd422: brom_out <= 64'd8621600869213436429;
    11'd423: brom_out <= 64'd2096562748759611565;
    11'd424: brom_out <= 64'd8349278891497519239;
    11'd425: brom_out <= 64'd346923801074208388;
    11'd426: brom_out <= 64'd6367974081209054997;
    11'd427: brom_out <= 64'd5762383813746039724;
    11'd428: brom_out <= 64'd1972299115398113399;
    11'd429: brom_out <= 64'd3713189838516711778;
    11'd430: brom_out <= 64'd1197769520636710353;
    11'd431: brom_out <= 64'd5608723318366677580;
    11'd432: brom_out <= 64'd3559594993567324157;
    11'd433: brom_out <= 64'd4575193000577835483;
    11'd434: brom_out <= 64'd3660689300204311631;
    11'd435: brom_out <= 64'd2416431477654523689;
    11'd436: brom_out <= 64'd4650911666456009623;
    11'd437: brom_out <= 64'd7522381762160574393;
    11'd438: brom_out <= 64'd190672817787439316;
    11'd439: brom_out <= 64'd325934885020391055;
    11'd440: brom_out <= 64'd706629558608325320;
    11'd441: brom_out <= 64'd3032300589071702614;
    11'd442: brom_out <= 64'd2579523930497909642;
    11'd443: brom_out <= 64'd2788024861033399442;
    11'd444: brom_out <= 64'd9002597627908969313;
    11'd445: brom_out <= 64'd6723624276537951429;
    11'd446: brom_out <= 64'd2608111876007635512;
    11'd447: brom_out <= 64'd2541081846948700755;
    11'd448: brom_out <= 64'd4659765458083320719;
    11'd449: brom_out <= 64'd3928376956683301646;
    11'd450: brom_out <= 64'd142053923599972979;
    11'd451: brom_out <= 64'd19360041183212556;
    11'd452: brom_out <= 64'd6857245434418581628;
    11'd453: brom_out <= 64'd2410203915673962172;
    11'd454: brom_out <= 64'd342621247588169017;
    11'd455: brom_out <= 64'd5315893553516886003;
    11'd456: brom_out <= 64'd7281806063522646650;
    11'd457: brom_out <= 64'd8410046497771752776;
    11'd458: brom_out <= 64'd2485207109882000355;
    11'd459: brom_out <= 64'd841862554873101340;
    11'd460: brom_out <= 64'd8519167899099856799;
    11'd461: brom_out <= 64'd4696904235291685297;
    11'd462: brom_out <= 64'd4270274588157767362;
    11'd463: brom_out <= 64'd7097500566651828779;
    11'd464: brom_out <= 64'd3865593938793959904;
    11'd465: brom_out <= 64'd4355722000643974519;
    11'd466: brom_out <= 64'd3970048001387779941;
    11'd467: brom_out <= 64'd1209619758992703366;
    11'd468: brom_out <= 64'd5514005748138490513;
    11'd469: brom_out <= 64'd688007168033240;
    11'd470: brom_out <= 64'd6999880349491995737;
    11'd471: brom_out <= 64'd4848939826616760681;
    11'd472: brom_out <= 64'd1198684013469568818;
    11'd473: brom_out <= 64'd8135295486259970094;
    11'd474: brom_out <= 64'd7830295104395985050;
    11'd475: brom_out <= 64'd7581053371999636081;
    11'd476: brom_out <= 64'd7931101422433936750;
    11'd477: brom_out <= 64'd2116647075839881756;
    11'd478: brom_out <= 64'd6703239196443292823;
    11'd479: brom_out <= 64'd7650526928209470539;
    11'd480: brom_out <= 64'd2401188481327814690;
    11'd481: brom_out <= 64'd850988766213502686;
    11'd482: brom_out <= 64'd2045199198493182244;
    11'd483: brom_out <= 64'd2618127369391731462;
    11'd484: brom_out <= 64'd7903854980513516255;
    11'd485: brom_out <= 64'd2094334658668413523;
    11'd486: brom_out <= 64'd2972592356844292403;
    11'd487: brom_out <= 64'd5176039432325527339;
    11'd488: brom_out <= 64'd4832896826743834449;
    11'd489: brom_out <= 64'd3820875116947407203;
    11'd490: brom_out <= 64'd4057810512372530111;
    11'd491: brom_out <= 64'd1830741857931679868;
    11'd492: brom_out <= 64'd7413850612596629259;
    11'd493: brom_out <= 64'd1797516723013854300;
    11'd494: brom_out <= 64'd5141180020896888574;
    11'd495: brom_out <= 64'd3777853455353424430;
    11'd496: brom_out <= 64'd2002943968299338895;
    11'd497: brom_out <= 64'd105518862569412047;
    11'd498: brom_out <= 64'd8659675561336273669;
    11'd499: brom_out <= 64'd4580270149773429686;
    11'd500: brom_out <= 64'd5789621183771780820;
    11'd501: brom_out <= 64'd3391235165647737720;
    11'd502: brom_out <= 64'd6400593500865891530;
    11'd503: brom_out <= 64'd3635580377175485895;
    11'd504: brom_out <= 64'd1406596659207299326;
    11'd505: brom_out <= 64'd3400202999108630343;
    11'd506: brom_out <= 64'd5039245648445919963;
    11'd507: brom_out <= 64'd6304614544456206336;
    11'd508: brom_out <= 64'd7546852068187909855;
    11'd509: brom_out <= 64'd4056535390267703032;
    11'd510: brom_out <= 64'd6049701732477573686;
    11'd511: brom_out <= 64'd7696362086031279642;
    11'd512: brom_out <= 64'd5694819423089841067;
    11'd513: brom_out <= 64'd8431301469303948298;
    11'd514: brom_out <= 64'd2413300624007091572;
    11'd515: brom_out <= 64'd3676771400266117330;
    11'd516: brom_out <= 64'd1439455466828941644;
    11'd517: brom_out <= 64'd2471528734300932856;
    11'd518: brom_out <= 64'd4935478512406328489;
    11'd519: brom_out <= 64'd4832653183844613201;
    11'd520: brom_out <= 64'd6991420717518923369;
    11'd521: brom_out <= 64'd4885623610012298224;
    11'd522: brom_out <= 64'd2698824602216536714;
    11'd523: brom_out <= 64'd4541017139054292672;
    11'd524: brom_out <= 64'd523263350017325961;
    11'd525: brom_out <= 64'd6200187860148334423;
    11'd526: brom_out <= 64'd2112942291044247589;
    11'd527: brom_out <= 64'd4741985617453118740;
    11'd528: brom_out <= 64'd3199971649867813866;
    11'd529: brom_out <= 64'd9199614664125632230;
    11'd530: brom_out <= 64'd721893744040243775;
    11'd531: brom_out <= 64'd6797302604172576659;
    11'd532: brom_out <= 64'd630226834235528396;
    11'd533: brom_out <= 64'd1288370651736466684;
    11'd534: brom_out <= 64'd6703339429733610384;
    11'd535: brom_out <= 64'd165369273176347238;
    11'd536: brom_out <= 64'd222948241930436619;
    11'd537: brom_out <= 64'd3625135611903007760;
    11'd538: brom_out <= 64'd6265219356917378798;
    11'd539: brom_out <= 64'd6212389645631186009;
    11'd540: brom_out <= 64'd2494091564964353659;
    11'd541: brom_out <= 64'd8746707750626208732;
    11'd542: brom_out <= 64'd9060509806960703546;
    11'd543: brom_out <= 64'd1464686228147214000;
    11'd544: brom_out <= 64'd2128614640918203358;
    11'd545: brom_out <= 64'd8226994774224310546;
    11'd546: brom_out <= 64'd2455922524235164580;
    11'd547: brom_out <= 64'd6421251889202531258;
    11'd548: brom_out <= 64'd5740686176908711475;
    11'd549: brom_out <= 64'd7839021458130261443;
    11'd550: brom_out <= 64'd3523071753482109712;
    11'd551: brom_out <= 64'd8999051484295950071;
    11'd552: brom_out <= 64'd6380027571086152967;
    11'd553: brom_out <= 64'd2582554806539286758;
    11'd554: brom_out <= 64'd7797469498989570118;
    11'd555: brom_out <= 64'd7149760397640115984;
    11'd556: brom_out <= 64'd5407165014541058846;
    11'd557: brom_out <= 64'd2488043764664355060;
    11'd558: brom_out <= 64'd3117944430576875629;
    11'd559: brom_out <= 64'd3932861293713858077;
    11'd560: brom_out <= 64'd4541486265004346961;
    11'd561: brom_out <= 64'd6508989279226413174;
    11'd562: brom_out <= 64'd143791927335086860;
    11'd563: brom_out <= 64'd1929632205213301446;
    11'd564: brom_out <= 64'd9161157683831349932;
    11'd565: brom_out <= 64'd2197388356117334702;
    11'd566: brom_out <= 64'd2691767668631111291;
    11'd567: brom_out <= 64'd3185863346693743704;
    11'd568: brom_out <= 64'd8930375953653963134;
    11'd569: brom_out <= 64'd7118858597288346597;
    11'd570: brom_out <= 64'd319884686633943643;
    11'd571: brom_out <= 64'd4323834995363520338;
    11'd572: brom_out <= 64'd2101313952790077927;
    11'd573: brom_out <= 64'd645892561257917929;
    11'd574: brom_out <= 64'd399969658011778878;
    11'd575: brom_out <= 64'd2598428332710975178;
    11'd576: brom_out <= 64'd7146228324775845589;
    11'd577: brom_out <= 64'd8631050930890094081;
    11'd578: brom_out <= 64'd7210109378417634812;
    11'd579: brom_out <= 64'd4014149304146885558;
    11'd580: brom_out <= 64'd7699005035771607412;
    11'd581: brom_out <= 64'd4449366486177894711;
    11'd582: brom_out <= 64'd3880882356684911754;
    11'd583: brom_out <= 64'd8458326417131546409;
    11'd584: brom_out <= 64'd2512504148219754733;
    11'd585: brom_out <= 64'd930503605682625418;
    11'd586: brom_out <= 64'd1171194988591484366;
    11'd587: brom_out <= 64'd915086647165685112;
    11'd588: brom_out <= 64'd6198596474422823906;
    11'd589: brom_out <= 64'd5213098489073531483;
    11'd590: brom_out <= 64'd1760832019471425278;
    11'd591: brom_out <= 64'd1538198027913715822;
    11'd592: brom_out <= 64'd1321928960272271311;
    11'd593: brom_out <= 64'd8029737381391845490;
    11'd594: brom_out <= 64'd2820343168317509442;
    11'd595: brom_out <= 64'd1214813679580018107;
    11'd596: brom_out <= 64'd5321756606589496737;
    11'd597: brom_out <= 64'd4217049811595050524;
    11'd598: brom_out <= 64'd3272746968595445449;
    11'd599: brom_out <= 64'd6335530199418981784;
    11'd600: brom_out <= 64'd2036924386199742561;
    11'd601: brom_out <= 64'd6674507905629246363;
    11'd602: brom_out <= 64'd7822652083037999802;
    11'd603: brom_out <= 64'd1421918644939809259;
    11'd604: brom_out <= 64'd608887493271275624;
    11'd605: brom_out <= 64'd6220940958186282004;
    11'd606: brom_out <= 64'd3674999362557584310;
    11'd607: brom_out <= 64'd8892259573730330161;
    11'd608: brom_out <= 64'd2620821568285243738;
    11'd609: brom_out <= 64'd6678854173437392197;
    11'd610: brom_out <= 64'd8954372130952231580;
    11'd611: brom_out <= 64'd8217059487227195162;
    11'd612: brom_out <= 64'd2756717500342111516;
    11'd613: brom_out <= 64'd8463007374782694281;
    11'd614: brom_out <= 64'd4905273512459903447;
    11'd615: brom_out <= 64'd5702571964487734279;
    11'd616: brom_out <= 64'd1745775350037015008;
    11'd617: brom_out <= 64'd5551820442000920135;
    11'd618: brom_out <= 64'd1045866548808442081;
    11'd619: brom_out <= 64'd2065426583040156382;
    11'd620: brom_out <= 64'd5349820788321212586;
    11'd621: brom_out <= 64'd514622884702815980;
    11'd622: brom_out <= 64'd761434371403642555;
    11'd623: brom_out <= 64'd4014438828781610649;
    11'd624: brom_out <= 64'd2645026052511064389;
    11'd625: brom_out <= 64'd5121860646049111138;
    11'd626: brom_out <= 64'd3433122314438944598;
    11'd627: brom_out <= 64'd8225186588976509856;
    11'd628: brom_out <= 64'd3543633365011365493;
    11'd629: brom_out <= 64'd9034265768767752860;
    11'd630: brom_out <= 64'd479232571601645093;
    11'd631: brom_out <= 64'd3956102820918726636;
    11'd632: brom_out <= 64'd1424284277694739202;
    11'd633: brom_out <= 64'd7115057179722603849;
    11'd634: brom_out <= 64'd8588788152872033952;
    11'd635: brom_out <= 64'd3299388022939274935;
    11'd636: brom_out <= 64'd3399641655016048048;
    11'd637: brom_out <= 64'd4215899052489957961;
    11'd638: brom_out <= 64'd3873611136974020819;
    11'd639: brom_out <= 64'd2051128225809906454;
    11'd640: brom_out <= 64'd4598343537641952316;
    11'd641: brom_out <= 64'd5430075770190133814;
    11'd642: brom_out <= 64'd8367401985994315753;
    11'd643: brom_out <= 64'd5780549035734671464;
    11'd644: brom_out <= 64'd6788515364259461350;
    11'd645: brom_out <= 64'd8126670364120682383;
    11'd646: brom_out <= 64'd5490110473127369071;
    11'd647: brom_out <= 64'd7019920813760977335;
    11'd648: brom_out <= 64'd1068506085308168299;
    11'd649: brom_out <= 64'd3160804074042342377;
    11'd650: brom_out <= 64'd4991872375415097966;
    11'd651: brom_out <= 64'd6748231796581112054;
    11'd652: brom_out <= 64'd535489186106420171;
    11'd653: brom_out <= 64'd3958739186601675842;
    11'd654: brom_out <= 64'd2675157303987172335;
    11'd655: brom_out <= 64'd797330655875880193;
    11'd656: brom_out <= 64'd6408137736931057484;
    11'd657: brom_out <= 64'd4850759160253046498;
    11'd658: brom_out <= 64'd6232318510873924032;
    11'd659: brom_out <= 64'd2599834517819486921;
    11'd660: brom_out <= 64'd5641334475235667248;
    11'd661: brom_out <= 64'd1203055569162238986;
    11'd662: brom_out <= 64'd5338323249244987111;
    11'd663: brom_out <= 64'd4247710559793395244;
    11'd664: brom_out <= 64'd8043843428201761120;
    11'd665: brom_out <= 64'd5199563489232049520;
    11'd666: brom_out <= 64'd2408995380763836064;
    11'd667: brom_out <= 64'd4007939317173556756;
    11'd668: brom_out <= 64'd2988003291163597772;
    11'd669: brom_out <= 64'd8527041029612690685;
    11'd670: brom_out <= 64'd5975042846443655256;
    11'd671: brom_out <= 64'd4154061164191240553;
    11'd672: brom_out <= 64'd6926649083160067776;
    11'd673: brom_out <= 64'd6959120323656798202;
    11'd674: brom_out <= 64'd3356085635373983500;
    11'd675: brom_out <= 64'd7450440303901916080;
    11'd676: brom_out <= 64'd4070759535854596369;
    11'd677: brom_out <= 64'd7590266728843860201;
    11'd678: brom_out <= 64'd7567059777563118840;
    11'd679: brom_out <= 64'd3997353415390603130;
    11'd680: brom_out <= 64'd2866365310898254699;
    11'd681: brom_out <= 64'd8018956454409193985;
    11'd682: brom_out <= 64'd281297336415387058;
    11'd683: brom_out <= 64'd5705449768401225063;
    11'd684: brom_out <= 64'd6954573009345611546;
    11'd685: brom_out <= 64'd2196134131328854202;
    11'd686: brom_out <= 64'd8963468084008150228;
    11'd687: brom_out <= 64'd4806833545128666290;
    11'd688: brom_out <= 64'd5856405985550173159;
    11'd689: brom_out <= 64'd6524060390258113390;
    11'd690: brom_out <= 64'd8684039960416699458;
    11'd691: brom_out <= 64'd6539381008209602217;
    11'd692: brom_out <= 64'd3984980496255740925;
    11'd693: brom_out <= 64'd5808747171359760037;
    11'd694: brom_out <= 64'd6820273228561734778;
    11'd695: brom_out <= 64'd4623445673059349627;
    11'd696: brom_out <= 64'd821122352901815804;
    11'd697: brom_out <= 64'd2297512628000869070;
    11'd698: brom_out <= 64'd259454704045312389;
    11'd699: brom_out <= 64'd4359908600724727113;
    11'd700: brom_out <= 64'd4165309535333037889;
    11'd701: brom_out <= 64'd8556724613961862630;
    11'd702: brom_out <= 64'd2443810846363983242;
    11'd703: brom_out <= 64'd5896557942093509657;
    11'd704: brom_out <= 64'd8724544381459047665;
    11'd705: brom_out <= 64'd2901923088602051584;
    11'd706: brom_out <= 64'd6746020898894390783;
    11'd707: brom_out <= 64'd6416881649853854070;
    11'd708: brom_out <= 64'd6734045381418689149;
    11'd709: brom_out <= 64'd8238511228338902902;
    11'd710: brom_out <= 64'd5707050340337892907;
    11'd711: brom_out <= 64'd2335661004110044355;
    11'd712: brom_out <= 64'd6700421300865381064;
    11'd713: brom_out <= 64'd8896743906568536409;
    11'd714: brom_out <= 64'd268149779945592459;
    11'd715: brom_out <= 64'd751586876332682772;
    11'd716: brom_out <= 64'd4225632203196813442;
    11'd717: brom_out <= 64'd6435187536035377203;
    11'd718: brom_out <= 64'd7644517197190347411;
    11'd719: brom_out <= 64'd1253063413056104552;
    11'd720: brom_out <= 64'd1009828133023932836;
    11'd721: brom_out <= 64'd6358448171523864630;
    11'd722: brom_out <= 64'd2015945304789420789;
    11'd723: brom_out <= 64'd695558424770826551;
    11'd724: brom_out <= 64'd4141171787133538854;
    11'd725: brom_out <= 64'd6252461585230888043;
    11'd726: brom_out <= 64'd4718646014166511125;
    11'd727: brom_out <= 64'd3995630726086934628;
    11'd728: brom_out <= 64'd1673544521435346038;
    11'd729: brom_out <= 64'd5183485982849115904;
    11'd730: brom_out <= 64'd3977574710926867577;
    11'd731: brom_out <= 64'd8883490896537391258;
    11'd732: brom_out <= 64'd268423085928125282;
    11'd733: brom_out <= 64'd2613352977137571904;
    11'd734: brom_out <= 64'd3172806986990922073;
    11'd735: brom_out <= 64'd673651761159149151;
    11'd736: brom_out <= 64'd2148959679869540120;
    11'd737: brom_out <= 64'd6762824372060873885;
    11'd738: brom_out <= 64'd8551686576092683850;
    11'd739: brom_out <= 64'd1007192545845825904;
    11'd740: brom_out <= 64'd3959612675003995092;
    11'd741: brom_out <= 64'd8738899863672466343;
    11'd742: brom_out <= 64'd4547765830837227036;
    11'd743: brom_out <= 64'd7119625349764498718;
    11'd744: brom_out <= 64'd3148100078089732519;
    11'd745: brom_out <= 64'd4246176443449053244;
    11'd746: brom_out <= 64'd6790481463797119064;
    11'd747: brom_out <= 64'd3449763520287903007;
    11'd748: brom_out <= 64'd3145191905961267984;
    11'd749: brom_out <= 64'd1905921935244999538;
    11'd750: brom_out <= 64'd3871541686777961704;
    11'd751: brom_out <= 64'd8729097820477921361;
    11'd752: brom_out <= 64'd5474825609301500618;
    11'd753: brom_out <= 64'd418407510091815277;
    11'd754: brom_out <= 64'd2764561907159231818;
    11'd755: brom_out <= 64'd6173199079945490225;
    11'd756: brom_out <= 64'd5335826789442547812;
    11'd757: brom_out <= 64'd5400690615858132495;
    11'd758: brom_out <= 64'd1501601289626383463;
    11'd759: brom_out <= 64'd4716183757898382283;
    11'd760: brom_out <= 64'd2400374672458484165;
    11'd761: brom_out <= 64'd6238947467064753318;
    11'd762: brom_out <= 64'd5328340207630532751;
    11'd763: brom_out <= 64'd98267416648275707;
    11'd764: brom_out <= 64'd4637045799031159911;
    11'd765: brom_out <= 64'd7906959063152076048;
    11'd766: brom_out <= 64'd7306985850419918102;
    11'd767: brom_out <= 64'd8891666758032158567;
    11'd768: brom_out <= 64'd4133337517863562233;
    11'd769: brom_out <= 64'd3027692497507765209;
    11'd770: brom_out <= 64'd7713485600285780027;
    11'd771: brom_out <= 64'd4171994359517618376;
    11'd772: brom_out <= 64'd9056522580924845506;
    11'd773: brom_out <= 64'd6895955466386430136;
    11'd774: brom_out <= 64'd5146944127070654897;
    11'd775: brom_out <= 64'd1536662417349835217;
    11'd776: brom_out <= 64'd7895346649673647512;
    11'd777: brom_out <= 64'd1615980629658654598;
    11'd778: brom_out <= 64'd6536782322229948227;
    11'd779: brom_out <= 64'd2604011659228572151;
    11'd780: brom_out <= 64'd6036498926837986101;
    11'd781: brom_out <= 64'd6441390040726608280;
    11'd782: brom_out <= 64'd3638521861921191001;
    11'd783: brom_out <= 64'd9000604085325519922;
    11'd784: brom_out <= 64'd2553480831479574171;
    11'd785: brom_out <= 64'd5605517858865043016;
    11'd786: brom_out <= 64'd9090913341983878540;
    11'd787: brom_out <= 64'd3354937147210049242;
    11'd788: brom_out <= 64'd8407678306248906235;
    11'd789: brom_out <= 64'd973208025566076311;
    11'd790: brom_out <= 64'd7410439247127875940;
    11'd791: brom_out <= 64'd6835377452905998223;
    11'd792: brom_out <= 64'd2154994274453286679;
    11'd793: brom_out <= 64'd3363071006717555626;
    11'd794: brom_out <= 64'd3411793274425605700;
    11'd795: brom_out <= 64'd643033505655820275;
    11'd796: brom_out <= 64'd186864364587700322;
    11'd797: brom_out <= 64'd3271882312209193996;
    11'd798: brom_out <= 64'd8201679816666974562;
    11'd799: brom_out <= 64'd6053585916959618025;
    11'd800: brom_out <= 64'd5338966768282452435;
    11'd801: brom_out <= 64'd8043406520314475049;
    11'd802: brom_out <= 64'd2217802334457014631;
    11'd803: brom_out <= 64'd3014029263312094735;
    11'd804: brom_out <= 64'd6583292799783687284;
    11'd805: brom_out <= 64'd3189914079696153009;
    11'd806: brom_out <= 64'd4138734928065873534;
    11'd807: brom_out <= 64'd4197947585696717855;
    11'd808: brom_out <= 64'd1482359963028216865;
    11'd809: brom_out <= 64'd8392599323902861453;
    11'd810: brom_out <= 64'd3076372057811423577;
    11'd811: brom_out <= 64'd3378640241265400310;
    11'd812: brom_out <= 64'd2530176121340192890;
    11'd813: brom_out <= 64'd6632009698444613753;
    11'd814: brom_out <= 64'd3422585145867265642;
    11'd815: brom_out <= 64'd3941604185467133427;
    11'd816: brom_out <= 64'd1352806655029681034;
    11'd817: brom_out <= 64'd7549902755199667399;
    11'd818: brom_out <= 64'd709496652131180917;
    11'd819: brom_out <= 64'd4117702578170040672;
    11'd820: brom_out <= 64'd8637989573606132378;
    11'd821: brom_out <= 64'd5807769899454577531;
    11'd822: brom_out <= 64'd354275588959183915;
    11'd823: brom_out <= 64'd296328949872700347;
    11'd824: brom_out <= 64'd3346591847539295845;
    11'd825: brom_out <= 64'd5281549017633074463;
    11'd826: brom_out <= 64'd2007220908801309791;
    11'd827: brom_out <= 64'd5349785661207910397;
    11'd828: brom_out <= 64'd2424397614063191733;
    11'd829: brom_out <= 64'd7222706162509528069;
    11'd830: brom_out <= 64'd1007320226254812508;
    11'd831: brom_out <= 64'd3018234359963511924;
    11'd832: brom_out <= 64'd7302840033919719354;
    11'd833: brom_out <= 64'd2968054662555921271;
    11'd834: brom_out <= 64'd8797336147399983457;
    11'd835: brom_out <= 64'd7077504767923673293;
    11'd836: brom_out <= 64'd3714939630179512644;
    11'd837: brom_out <= 64'd3847814091255260418;
    11'd838: brom_out <= 64'd291704881778621267;
    11'd839: brom_out <= 64'd1890046659933707987;
    11'd840: brom_out <= 64'd4657523443218805420;
    11'd841: brom_out <= 64'd7289874174738232147;
    11'd842: brom_out <= 64'd5261056114704450048;
    11'd843: brom_out <= 64'd6075870574138795397;
    11'd844: brom_out <= 64'd44734367532455404;
    11'd845: brom_out <= 64'd120845593022123278;
    11'd846: brom_out <= 64'd8461716466987517362;
    11'd847: brom_out <= 64'd7365794054744162278;
    11'd848: brom_out <= 64'd2700680744585487300;
    11'd849: brom_out <= 64'd370793600216804065;
    11'd850: brom_out <= 64'd1777888570579566155;
    11'd851: brom_out <= 64'd6620688383163974071;
    11'd852: brom_out <= 64'd203579238871197068;
    11'd853: brom_out <= 64'd1638450655490297613;
    11'd854: brom_out <= 64'd7029508759137299187;
    11'd855: brom_out <= 64'd8894609215971099829;
    11'd856: brom_out <= 64'd824780095341126479;
    11'd857: brom_out <= 64'd7854543062470227875;
    11'd858: brom_out <= 64'd8629464100960320937;
    11'd859: brom_out <= 64'd5449865088360881617;
    11'd860: brom_out <= 64'd4194926527731236764;
    11'd861: brom_out <= 64'd2039700583643793626;
    11'd862: brom_out <= 64'd7666856413403412022;
    11'd863: brom_out <= 64'd5445771681671222660;
    11'd864: brom_out <= 64'd4441256879323813867;
    11'd865: brom_out <= 64'd4371251341607182761;
    11'd866: brom_out <= 64'd8599591383127997894;
    11'd867: brom_out <= 64'd4347545940856227957;
    11'd868: brom_out <= 64'd989263098681289775;
    11'd869: brom_out <= 64'd7064390324490644869;
    11'd870: brom_out <= 64'd6120494681119218490;
    11'd871: brom_out <= 64'd6307135453118974578;
    11'd872: brom_out <= 64'd8320486820135076887;
    11'd873: brom_out <= 64'd2053859704017476493;
    11'd874: brom_out <= 64'd1805999465650818267;
    11'd875: brom_out <= 64'd5123132371367846493;
    11'd876: brom_out <= 64'd8506952230442773713;
    11'd877: brom_out <= 64'd6174441468423999837;
    11'd878: brom_out <= 64'd6952577279346250668;
    11'd879: brom_out <= 64'd8404272663876270125;
    11'd880: brom_out <= 64'd7142821866876178327;
    11'd881: brom_out <= 64'd8720908108610768275;
    11'd882: brom_out <= 64'd2656869541187597167;
    11'd883: brom_out <= 64'd7535490219096512345;
    11'd884: brom_out <= 64'd3431191520018159239;
    11'd885: brom_out <= 64'd7910040705147176291;
    11'd886: brom_out <= 64'd7349482934862272877;
    11'd887: brom_out <= 64'd7597426467432823857;
    11'd888: brom_out <= 64'd1481948738260612947;
    11'd889: brom_out <= 64'd8821216360349768285;
    11'd890: brom_out <= 64'd6912811304509913612;
    11'd891: brom_out <= 64'd1919407470247348674;
    11'd892: brom_out <= 64'd7059253706224036243;
    11'd893: brom_out <= 64'd8597923735828669071;
    11'd894: brom_out <= 64'd7285101071736128928;
    11'd895: brom_out <= 64'd3555685980750069891;
    11'd896: brom_out <= 64'd3423547344888630074;
    11'd897: brom_out <= 64'd2233404176129745739;
    11'd898: brom_out <= 64'd5516120319229414306;
    11'd899: brom_out <= 64'd7085601456569950070;
    11'd900: brom_out <= 64'd7330712937655359649;
    11'd901: brom_out <= 64'd172307991973364026;
    11'd902: brom_out <= 64'd3674227907828554084;
    11'd903: brom_out <= 64'd2119460563244100556;
    11'd904: brom_out <= 64'd9108416585855612745;
    11'd905: brom_out <= 64'd3326407409724130966;
    11'd906: brom_out <= 64'd8260964555008341506;
    11'd907: brom_out <= 64'd7871198280510774602;
    11'd908: brom_out <= 64'd7478335139546753414;
    11'd909: brom_out <= 64'd4179314389048712511;
    11'd910: brom_out <= 64'd7017007038818110112;
    11'd911: brom_out <= 64'd8769561004090428205;
    11'd912: brom_out <= 64'd806930591695923861;
    11'd913: brom_out <= 64'd8140052029682996333;
    11'd914: brom_out <= 64'd7909088071210934417;
    11'd915: brom_out <= 64'd3484417785571238429;
    11'd916: brom_out <= 64'd4051896663704402160;
    11'd917: brom_out <= 64'd1563022718788315335;
    11'd918: brom_out <= 64'd3964592748051227703;
    11'd919: brom_out <= 64'd2790516225524970165;
    11'd920: brom_out <= 64'd1385279684519564741;
    11'd921: brom_out <= 64'd3529697055032030879;
    11'd922: brom_out <= 64'd1067989342997180519;
    11'd923: brom_out <= 64'd235349974241710564;
    11'd924: brom_out <= 64'd3900620095247252000;
    11'd925: brom_out <= 64'd4445499959798319734;
    11'd926: brom_out <= 64'd6061538969494844847;
    11'd927: brom_out <= 64'd5383589726029507980;
    11'd928: brom_out <= 64'd8804992667951521152;
    11'd929: brom_out <= 64'd5140936975578878114;
    11'd930: brom_out <= 64'd1530938870927555532;
    11'd931: brom_out <= 64'd6791361877209584700;
    11'd932: brom_out <= 64'd1193864816184446735;
    11'd933: brom_out <= 64'd1617401520512653107;
    11'd934: brom_out <= 64'd5722470941604677021;
    11'd935: brom_out <= 64'd5322375988547217422;
    11'd936: brom_out <= 64'd3268957955472527918;
    11'd937: brom_out <= 64'd4421054392861095009;
    11'd938: brom_out <= 64'd2211632914135038092;
    11'd939: brom_out <= 64'd7891747589757095064;
    11'd940: brom_out <= 64'd2707564795335828269;
    11'd941: brom_out <= 64'd848659378860328351;
    11'd942: brom_out <= 64'd4084398432585418431;
    11'd943: brom_out <= 64'd1374371692087762288;
    11'd944: brom_out <= 64'd1309332277140087809;
    11'd945: brom_out <= 64'd6039700011317030473;
    11'd946: brom_out <= 64'd62208054836922472;
    11'd947: brom_out <= 64'd1975259188211765586;
    11'd948: brom_out <= 64'd5829687652731346729;
    11'd949: brom_out <= 64'd1552859820987002409;
    11'd950: brom_out <= 64'd4337357512006263771;
    11'd951: brom_out <= 64'd8804683524608505769;
    11'd952: brom_out <= 64'd1544044049239432418;
    11'd953: brom_out <= 64'd9198233257987748235;
    11'd954: brom_out <= 64'd325508699914523933;
    11'd955: brom_out <= 64'd7444143362807642230;
    11'd956: brom_out <= 64'd1301211514226427325;
    11'd957: brom_out <= 64'd7050308007514871294;
    11'd958: brom_out <= 64'd9058697836308692493;
    11'd959: brom_out <= 64'd1898187455399378490;
    11'd960: brom_out <= 64'd4425969977592900653;
    11'd961: brom_out <= 64'd5211508916412346537;
    11'd962: brom_out <= 64'd7337507285800242744;
    11'd963: brom_out <= 64'd8102267769625153817;
    11'd964: brom_out <= 64'd4374120169651761055;
    11'd965: brom_out <= 64'd5443168134129117719;
    11'd966: brom_out <= 64'd3018287891620215876;
    11'd967: brom_out <= 64'd1722440177768065768;
    11'd968: brom_out <= 64'd5692414573629404816;
    11'd969: brom_out <= 64'd291047870053758273;
    11'd970: brom_out <= 64'd5710927416131961609;
    11'd971: brom_out <= 64'd5395679680946821168;
    11'd972: brom_out <= 64'd123993695763643615;
    11'd973: brom_out <= 64'd2626948377526316580;
    11'd974: brom_out <= 64'd2927196191119788241;
    11'd975: brom_out <= 64'd4062878447447081317;
    11'd976: brom_out <= 64'd2961872907626903907;
    11'd977: brom_out <= 64'd5199136735088625411;
    11'd978: brom_out <= 64'd5459877254919301330;
    11'd979: brom_out <= 64'd5007789230245417606;
    11'd980: brom_out <= 64'd3007686203960454990;
    11'd981: brom_out <= 64'd8745252878040690631;
    11'd982: brom_out <= 64'd392878258471787806;
    11'd983: brom_out <= 64'd3278352673360321384;
    11'd984: brom_out <= 64'd8318291207326965041;
    11'd985: brom_out <= 64'd3061302262506944119;
    11'd986: brom_out <= 64'd4876711006616769883;
    11'd987: brom_out <= 64'd4809336419563746839;
    11'd988: brom_out <= 64'd5834673946691031217;
    11'd989: brom_out <= 64'd8888021460029350015;
    11'd990: brom_out <= 64'd4005169494037905846;
    11'd991: brom_out <= 64'd8878823148073529111;
    11'd992: brom_out <= 64'd4659246901878184726;
    11'd993: brom_out <= 64'd2000836378318539205;
    11'd994: brom_out <= 64'd2889893669248460690;
    11'd995: brom_out <= 64'd8019432184343326435;
    11'd996: brom_out <= 64'd2823155742120844428;
    11'd997: brom_out <= 64'd4310852202031595690;
    11'd998: brom_out <= 64'd2958226008256126502;
    11'd999: brom_out <= 64'd8033699588279788769;
    11'd1000: brom_out <= 64'd93431844872797265;
    11'd1001: brom_out <= 64'd5272789992716447134;
    11'd1002: brom_out <= 64'd1164853792565412535;
    11'd1003: brom_out <= 64'd4853549291935722968;
    11'd1004: brom_out <= 64'd3264067940062730346;
    11'd1005: brom_out <= 64'd7930951055937939494;
    11'd1006: brom_out <= 64'd822406158089873071;
    11'd1007: brom_out <= 64'd5520853189671187665;
    11'd1008: brom_out <= 64'd5306051938089152367;
    11'd1009: brom_out <= 64'd7709314815903447805;
    11'd1010: brom_out <= 64'd406871917756752571;
    11'd1011: brom_out <= 64'd1648603819215645742;
    11'd1012: brom_out <= 64'd5109171197189782695;
    11'd1013: brom_out <= 64'd5589392136524859205;
    11'd1014: brom_out <= 64'd1161635928050851819;
    11'd1015: brom_out <= 64'd7184851511033041049;
    11'd1016: brom_out <= 64'd9160988738586692345;
    11'd1017: brom_out <= 64'd9144850910909373196;
    11'd1018: brom_out <= 64'd5967134563948484553;
    11'd1019: brom_out <= 64'd6421505013862266551;
    11'd1020: brom_out <= 64'd6545306907600364841;
    11'd1021: brom_out <= 64'd5218254320364951087;
    11'd1022: brom_out <= 64'd4627640233359996770;
    11'd1023: brom_out <= 64'd8120458936301571092;
    default: brom_out <= 64'h1;
    endcase
end

generate
    if(DELAY == 1) begin
        assign b = brom_out;
    end
endgenerate

endmodule

//-------------------------------------------------------------------------------------------------

module tw_rom_11_intt_nwc
#(
    parameter LOGN  = 11,
    parameter LOGQ  = 64,
    parameter DELAY = 1,
    parameter STAGE = 11
)(
    input            clk,
    input [LOGN-1:0] raddr,
    output[LOGQ-1:0] b
);

(* ram_style = "block" *)
reg [LOGQ-1:0] brom_out, brom_out2;

always @(posedge clk) begin
    case(raddr[STAGE-1:0])
    12'd0: brom_out <= 64'd4800325891501495425;
    12'd1: brom_out <= 64'd3479955663905624912;
    12'd2: brom_out <= 64'd6942686573313721449;
    12'd3: brom_out <= 64'd2859865282093209065;
    12'd4: brom_out <= 64'd5499182698979939570;
    12'd5: brom_out <= 64'd2855896583733398539;
    12'd6: brom_out <= 64'd9195430145952975242;
    12'd7: brom_out <= 64'd268523678609812267;
    12'd8: brom_out <= 64'd3300993837355370774;
    12'd9: brom_out <= 64'd5779659341364002408;
    12'd10: brom_out <= 64'd6895474870082812174;
    12'd11: brom_out <= 64'd5417860397405817535;
    12'd12: brom_out <= 64'd3763063295663263880;
    12'd13: brom_out <= 64'd2035072135929394071;
    12'd14: brom_out <= 64'd8411697026915987727;
    12'd15: brom_out <= 64'd4207477549930981961;
    12'd16: brom_out <= 64'd2371121004762206413;
    12'd17: brom_out <= 64'd772015388505701109;
    12'd18: brom_out <= 64'd1291769418475865586;
    12'd19: brom_out <= 64'd9141993189948588563;
    12'd20: brom_out <= 64'd2162936514908913563;
    12'd21: brom_out <= 64'd1898016065535012275;
    12'd22: brom_out <= 64'd2528879447085842517;
    12'd23: brom_out <= 64'd2311408450510800010;
    12'd24: brom_out <= 64'd7507303259201390021;
    12'd25: brom_out <= 64'd4762074383448690520;
    12'd26: brom_out <= 64'd249568661117497673;
    12'd27: brom_out <= 64'd1518691922593280722;
    12'd28: brom_out <= 64'd659317911363937817;
    12'd29: brom_out <= 64'd3128431811455045720;
    12'd30: brom_out <= 64'd6190591306936762157;
    12'd31: brom_out <= 64'd2034678932731682912;
    12'd32: brom_out <= 64'd3077267012251774723;
    12'd33: brom_out <= 64'd5701780488963733939;
    12'd34: brom_out <= 64'd2691484975942555879;
    12'd35: brom_out <= 64'd526419352956882135;
    12'd36: brom_out <= 64'd3222150524692787156;
    12'd37: brom_out <= 64'd7264146735115973951;
    12'd38: brom_out <= 64'd398573074911215638;
    12'd39: brom_out <= 64'd8145476396298478751;
    12'd40: brom_out <= 64'd2505141805715690065;
    12'd41: brom_out <= 64'd4148880509067847681;
    12'd42: brom_out <= 64'd1316642780790498741;
    12'd43: brom_out <= 64'd6989158732632716781;
    12'd44: brom_out <= 64'd2851678937043902667;
    12'd45: brom_out <= 64'd6709388255283723070;
    12'd46: brom_out <= 64'd7816234934658379448;
    12'd47: brom_out <= 64'd4666785398365578624;
    12'd48: brom_out <= 64'd7934631291163394022;
    12'd49: brom_out <= 64'd1159284894254976374;
    12'd50: brom_out <= 64'd4243273064418189329;
    12'd51: brom_out <= 64'd3981921757822415978;
    12'd52: brom_out <= 64'd6691909628951155125;
    12'd53: brom_out <= 64'd2338193104926316584;
    12'd54: brom_out <= 64'd1663073629993296632;
    12'd55: brom_out <= 64'd7023774353635676184;
    12'd56: brom_out <= 64'd3378677374409253768;
    12'd57: brom_out <= 64'd6394875299066583771;
    12'd58: brom_out <= 64'd2374307618530860008;
    12'd59: brom_out <= 64'd5943036323825889194;
    12'd60: brom_out <= 64'd7613523031203569219;
    12'd61: brom_out <= 64'd6687702232866970904;
    12'd62: brom_out <= 64'd4053328842517216816;
    12'd63: brom_out <= 64'd4709098501258011541;
    12'd64: brom_out <= 64'd2374694900661844296;
    12'd65: brom_out <= 64'd1618288916964425384;
    12'd66: brom_out <= 64'd2772437297514657011;
    12'd67: brom_out <= 64'd5270785824266435531;
    12'd68: brom_out <= 64'd2396521636741935089;
    12'd69: brom_out <= 64'd4522583066803542678;
    12'd70: brom_out <= 64'd1058894820381756984;
    12'd71: brom_out <= 64'd8103776501554795239;
    12'd72: brom_out <= 64'd1257205976697436021;
    12'd73: brom_out <= 64'd2097906600216330458;
    12'd74: brom_out <= 64'd6286024435479652455;
    12'd75: brom_out <= 64'd2233217965831104691;
    12'd76: brom_out <= 64'd2941897417371093549;
    12'd77: brom_out <= 64'd4060143600394135002;
    12'd78: brom_out <= 64'd678912652673726946;
    12'd79: brom_out <= 64'd8395280712977132829;
    12'd80: brom_out <= 64'd7125284802318235209;
    12'd81: brom_out <= 64'd7558182034901277051;
    12'd82: brom_out <= 64'd1690394721022924538;
    12'd83: brom_out <= 64'd5412118970273754969;
    12'd84: brom_out <= 64'd5236825456431198728;
    12'd85: brom_out <= 64'd5395111291698076598;
    12'd86: brom_out <= 64'd6145624954448652370;
    12'd87: brom_out <= 64'd4407679216896856922;
    12'd88: brom_out <= 64'd6861048754277304935;
    12'd89: brom_out <= 64'd5157703172826989787;
    12'd90: brom_out <= 64'd8027685862106484926;
    12'd91: brom_out <= 64'd6802831625721368331;
    12'd92: brom_out <= 64'd2785053808996448559;
    12'd93: brom_out <= 64'd1991486632246496547;
    12'd94: brom_out <= 64'd8742269389515150308;
    12'd95: brom_out <= 64'd1862212185359501624;
    12'd96: brom_out <= 64'd6479389135574218089;
    12'd97: brom_out <= 64'd5797796918016986849;
    12'd98: brom_out <= 64'd8062420006207593658;
    12'd99: brom_out <= 64'd3957775192915183035;
    12'd100: brom_out <= 64'd4634701814857146924;
    12'd101: brom_out <= 64'd8725412177447277056;
    12'd102: brom_out <= 64'd4018650761969710447;
    12'd103: brom_out <= 64'd7292324541740260853;
    12'd104: brom_out <= 64'd849943903253009125;
    12'd105: brom_out <= 64'd431075052699718718;
    12'd106: brom_out <= 64'd7974987193888671641;
    12'd107: brom_out <= 64'd712922527871334585;
    12'd108: brom_out <= 64'd3800294078297268779;
    12'd109: brom_out <= 64'd8095584328242765021;
    12'd110: brom_out <= 64'd9089338015047633280;
    12'd111: brom_out <= 64'd5601327057638316266;
    12'd112: brom_out <= 64'd8649892222598786589;
    12'd113: brom_out <= 64'd3210270500191530901;
    12'd114: brom_out <= 64'd5151280726591025649;
    12'd115: brom_out <= 64'd7147556857556972914;
    12'd116: brom_out <= 64'd7766075252890350202;
    12'd117: brom_out <= 64'd5480464217302446705;
    12'd118: brom_out <= 64'd6476766801164997754;
    12'd119: brom_out <= 64'd2597273667992680221;
    12'd120: brom_out <= 64'd3790452324141925863;
    12'd121: brom_out <= 64'd4794040938066575215;
    12'd122: brom_out <= 64'd2589582939823414234;
    12'd123: brom_out <= 64'd756466048455930835;
    12'd124: brom_out <= 64'd2966549754675922566;
    12'd125: brom_out <= 64'd6226886595030389768;
    12'd126: brom_out <= 64'd1496660390337478612;
    12'd127: brom_out <= 64'd6657664286413801039;
    12'd128: brom_out <= 64'd6222745039014399876;
    12'd129: brom_out <= 64'd426301473220411395;
    12'd130: brom_out <= 64'd4859005696659248678;
    12'd131: brom_out <= 64'd3630644555464587741;
    12'd132: brom_out <= 64'd2416324748724178781;
    12'd133: brom_out <= 64'd1236969277230738101;
    12'd134: brom_out <= 64'd377097061317563800;
    12'd135: brom_out <= 64'd2159646420240227088;
    12'd136: brom_out <= 64'd8512893223122605373;
    12'd137: brom_out <= 64'd4819778497996814306;
    12'd138: brom_out <= 64'd1537523827651003953;
    12'd139: brom_out <= 64'd3439788089689583316;
    12'd140: brom_out <= 64'd4316362393121156796;
    12'd141: brom_out <= 64'd4220445291959946550;
    12'd142: brom_out <= 64'd1910565994514953738;
    12'd143: brom_out <= 64'd3386790625943016997;
    12'd144: brom_out <= 64'd259562526787940444;
    12'd145: brom_out <= 64'd2299243199755714738;
    12'd146: brom_out <= 64'd6986793039503755230;
    12'd147: brom_out <= 64'd1511973552337218705;
    12'd148: brom_out <= 64'd4562119421056321697;
    12'd149: brom_out <= 64'd3239732047188120862;
    12'd150: brom_out <= 64'd7697589950031188899;
    12'd151: brom_out <= 64'd1018695198542940947;
    12'd152: brom_out <= 64'd3252396083063158562;
    12'd153: brom_out <= 64'd1241392538994811678;
    12'd154: brom_out <= 64'd2530669113643804885;
    12'd155: brom_out <= 64'd212665923330336927;
    12'd156: brom_out <= 64'd665408824541600341;
    12'd157: brom_out <= 64'd6791904410913986857;
    12'd158: brom_out <= 64'd7721772775943974989;
    12'd159: brom_out <= 64'd5055521811016418548;
    12'd160: brom_out <= 64'd3452367604655046608;
    12'd161: brom_out <= 64'd4750671555136292390;
    12'd162: brom_out <= 64'd6969456975579668172;
    12'd163: brom_out <= 64'd661923266498850602;
    12'd164: brom_out <= 64'd541897457463837983;
    12'd165: brom_out <= 64'd2701646318137365251;
    12'd166: brom_out <= 64'd1722905024214037943;
    12'd167: brom_out <= 64'd3670769217368925179;
    12'd168: brom_out <= 64'd7932816493105831575;
    12'd169: brom_out <= 64'd8850531379736829538;
    12'd170: brom_out <= 64'd7888051197376901843;
    12'd171: brom_out <= 64'd3425577606761650241;
    12'd172: brom_out <= 64'd1179206226387385431;
    12'd173: brom_out <= 64'd456151376233940003;
    12'd174: brom_out <= 64'd2156880501834892587;
    12'd175: brom_out <= 64'd6668291387187356098;
    12'd176: brom_out <= 64'd8133935149399888812;
    12'd177: brom_out <= 64'd1774899703521283622;
    12'd178: brom_out <= 64'd5875867150314008782;
    12'd179: brom_out <= 64'd5164053181159552141;
    12'd180: brom_out <= 64'd1713332285587794028;
    12'd181: brom_out <= 64'd7951951361044297533;
    12'd182: brom_out <= 64'd8146181411589677771;
    12'd183: brom_out <= 64'd6953870572822020170;
    12'd184: brom_out <= 64'd9196931934858870131;
    12'd185: brom_out <= 64'd5598363430607474864;
    12'd186: brom_out <= 64'd4648998823029332422;
    12'd187: brom_out <= 64'd700020304646857314;
    12'd188: brom_out <= 64'd5523662497685535193;
    12'd189: brom_out <= 64'd5152845739689556948;
    12'd190: brom_out <= 64'd7359435094937928283;
    12'd191: brom_out <= 64'd1125545921381746443;
    12'd192: brom_out <= 64'd2538395582094999318;
    12'd193: brom_out <= 64'd423630526441374453;
    12'd194: brom_out <= 64'd1820754629513803801;
    12'd195: brom_out <= 64'd1845376210427078657;
    12'd196: brom_out <= 64'd7368678072715404102;
    12'd197: brom_out <= 64'd7072358367783034174;
    12'd198: brom_out <= 64'd4162776424936148707;
    12'd199: brom_out <= 64'd7759374948081196863;
    12'd200: brom_out <= 64'd3010709835068914341;
    12'd201: brom_out <= 64'd3646902721873295276;
    12'd202: brom_out <= 64'd1147728471066900272;
    12'd203: brom_out <= 64'd7656339839612772097;
    12'd204: brom_out <= 64'd6054990505757038250;
    12'd205: brom_out <= 64'd1013679152589519969;
    12'd206: brom_out <= 64'd8333743826310743340;
    12'd207: brom_out <= 64'd3642594086284002188;
    12'd208: brom_out <= 64'd8500114950055893575;
    12'd209: brom_out <= 64'd3679758911276399796;
    12'd210: brom_out <= 64'd1783638055775460814;
    12'd211: brom_out <= 64'd8747729877227536812;
    12'd212: brom_out <= 64'd4329377037132016548;
    12'd213: brom_out <= 64'd3168697732681573307;
    12'd214: brom_out <= 64'd4206548617478432447;
    12'd215: brom_out <= 64'd464895284687076203;
    12'd216: brom_out <= 64'd8076401025279924364;
    12'd217: brom_out <= 64'd5267458570641341886;
    12'd218: brom_out <= 64'd8276971889301839992;
    12'd219: brom_out <= 64'd5898817955455751241;
    12'd220: brom_out <= 64'd698307562786839200;
    12'd221: brom_out <= 64'd5709904708196673668;
    12'd222: brom_out <= 64'd5241582045101281478;
    12'd223: brom_out <= 64'd9025568243707556001;
    12'd224: brom_out <= 64'd3055459869261096559;
    12'd225: brom_out <= 64'd5340937562885825391;
    12'd226: brom_out <= 64'd8194299551051940030;
    12'd227: brom_out <= 64'd3493583037585086015;
    12'd228: brom_out <= 64'd5356311159666381783;
    12'd229: brom_out <= 64'd3629269169643201619;
    12'd230: brom_out <= 64'd4524420868300376971;
    12'd231: brom_out <= 64'd6759275879853206024;
    12'd232: brom_out <= 64'd8552326562371205351;
    12'd233: brom_out <= 64'd7040166696894905205;
    12'd234: brom_out <= 64'd8217389348989696376;
    12'd235: brom_out <= 64'd4429484931225059437;
    12'd236: brom_out <= 64'd1641165469903478691;
    12'd237: brom_out <= 64'd1202078975675922520;
    12'd238: brom_out <= 64'd7959860158056540716;
    12'd239: brom_out <= 64'd2225169134372382396;
    12'd240: brom_out <= 64'd3227966121575495289;
    12'd241: brom_out <= 64'd7346350426691758711;
    12'd242: brom_out <= 64'd7020647700008759981;
    12'd243: brom_out <= 64'd5031825498998110876;
    12'd244: brom_out <= 64'd8199195365829297059;
    12'd245: brom_out <= 64'd7413771439580747971;
    12'd246: brom_out <= 64'd3139857114490429865;
    12'd247: brom_out <= 64'd8043870031834710239;
    12'd248: brom_out <= 64'd3778758662330671509;
    12'd249: brom_out <= 64'd8540671389212035800;
    12'd250: brom_out <= 64'd7902413825471882168;
    12'd251: brom_out <= 64'd5003737266267378347;
    12'd252: brom_out <= 64'd4222671849907000218;
    12'd253: brom_out <= 64'd4814619341200892449;
    12'd254: brom_out <= 64'd5731590892918121185;
    12'd255: brom_out <= 64'd8026654363533533980;
    12'd256: brom_out <= 64'd8896426049497849627;
    12'd257: brom_out <= 64'd6199835901485982447;
    12'd258: brom_out <= 64'd4376402107651772548;
    12'd259: brom_out <= 64'd2253757488076581512;
    12'd260: brom_out <= 64'd3093388195924954419;
    12'd261: brom_out <= 64'd1428513325448730781;
    12'd262: brom_out <= 64'd1504867771174291973;
    12'd263: brom_out <= 64'd5677691476163543173;
    12'd264: brom_out <= 64'd2391438443701480191;
    12'd265: brom_out <= 64'd695946579015900153;
    12'd266: brom_out <= 64'd7294996205506811847;
    12'd267: brom_out <= 64'd7988038772633490625;
    12'd268: brom_out <= 64'd2025129515112607752;
    12'd269: brom_out <= 64'd9191246919904120884;
    12'd270: brom_out <= 64'd859535790990336463;
    12'd271: brom_out <= 64'd4207798226736684758;
    12'd272: brom_out <= 64'd6688030206191899257;
    12'd273: brom_out <= 64'd2277697486818983507;
    12'd274: brom_out <= 64'd844050170434595647;
    12'd275: brom_out <= 64'd1490764820867971186;
    12'd276: brom_out <= 64'd627701391894460943;
    12'd277: brom_out <= 64'd2534636846613195505;
    12'd278: brom_out <= 64'd780097985034638355;
    12'd279: brom_out <= 64'd1749618515824061104;
    12'd280: brom_out <= 64'd5966825310262623229;
    12'd281: brom_out <= 64'd1453210662793346909;
    12'd282: brom_out <= 64'd7366540421523776714;
    12'd283: brom_out <= 64'd2420077835528011390;
    12'd284: brom_out <= 64'd495583132590109196;
    12'd285: brom_out <= 64'd6932768688618351052;
    12'd286: brom_out <= 64'd6551696432311407014;
    12'd287: brom_out <= 64'd6134086625494614808;
    12'd288: brom_out <= 64'd5366550186008764116;
    12'd289: brom_out <= 64'd4110532040090786872;
    12'd290: brom_out <= 64'd790096917042549410;
    12'd291: brom_out <= 64'd5541191997131717403;
    12'd292: brom_out <= 64'd3999844389222340392;
    12'd293: brom_out <= 64'd4120943426844979160;
    12'd294: brom_out <= 64'd7428861236385220425;
    12'd295: brom_out <= 64'd6639951088105649209;
    12'd296: brom_out <= 64'd2403990246273367937;
    12'd297: brom_out <= 64'd7447281614795883653;
    12'd298: brom_out <= 64'd7897746628230077827;
    12'd299: brom_out <= 64'd9149654981310430708;
    12'd300: brom_out <= 64'd3574747214061382244;
    12'd301: brom_out <= 64'd4749897991621604173;
    12'd302: brom_out <= 64'd8617949205266935393;
    12'd303: brom_out <= 64'd8121774868912873261;
    12'd304: brom_out <= 64'd2323165427717129126;
    12'd305: brom_out <= 64'd4083588380895555261;
    12'd306: brom_out <= 64'd8035095571273705487;
    12'd307: brom_out <= 64'd8493561211935137304;
    12'd308: brom_out <= 64'd8504628543831529531;
    12'd309: brom_out <= 64'd2436502221107518872;
    12'd310: brom_out <= 64'd5598789769912105197;
    12'd311: brom_out <= 64'd6489129592287459196;
    12'd312: brom_out <= 64'd7465755558447636714;
    12'd313: brom_out <= 64'd4657188657137503639;
    12'd314: brom_out <= 64'd182241072216388829;
    12'd315: brom_out <= 64'd5100059702679082872;
    12'd316: brom_out <= 64'd6692785604325659625;
    12'd317: brom_out <= 64'd2801845708307735242;
    12'd318: brom_out <= 64'd5491017919115305135;
    12'd319: brom_out <= 64'd9002871762156300039;
    12'd320: brom_out <= 64'd2149536796278676308;
    12'd321: brom_out <= 64'd3010964216135620168;
    12'd322: brom_out <= 64'd6781532021778605219;
    12'd323: brom_out <= 64'd4603521168701892011;
    12'd324: brom_out <= 64'd1833448269704610266;
    12'd325: brom_out <= 64'd1314124759094827101;
    12'd326: brom_out <= 64'd1151136055862584706;
    12'd327: brom_out <= 64'd8480587392932362214;
    12'd328: brom_out <= 64'd5936261658022389367;
    12'd329: brom_out <= 64'd7142156318395761314;
    12'd330: brom_out <= 64'd7762537989895041471;
    12'd331: brom_out <= 64'd6373218047476906700;
    12'd332: brom_out <= 64'd5729532631005382038;
    12'd333: brom_out <= 64'd2627914157997921697;
    12'd334: brom_out <= 64'd44571010367109978;
    12'd335: brom_out <= 64'd582202087413158924;
    12'd336: brom_out <= 64'd6382022418387363169;
    12'd337: brom_out <= 64'd5592765730425286444;
    12'd338: brom_out <= 64'd994769519486452848;
    12'd339: brom_out <= 64'd8862887296795875047;
    12'd340: brom_out <= 64'd8529148174397921760;
    12'd341: brom_out <= 64'd6869970591854709169;
    12'd342: brom_out <= 64'd3290498720694881330;
    12'd343: brom_out <= 64'd5646243182744253262;
    12'd344: brom_out <= 64'd7402905527746317978;
    12'd345: brom_out <= 64'd7370407779674085494;
    12'd346: brom_out <= 64'd3801989492430001416;
    12'd347: brom_out <= 64'd8432500509309037595;
    12'd348: brom_out <= 64'd1296704492479940580;
    12'd349: brom_out <= 64'd8542847765153714010;
    12'd350: brom_out <= 64'd3446805570613934959;
    12'd351: brom_out <= 64'd4305197521463115295;
    12'd352: brom_out <= 64'd8723174160948242557;
    12'd353: brom_out <= 64'd6685306183820187534;
    12'd354: brom_out <= 64'd4388567976140890533;
    12'd355: brom_out <= 64'd7748340154365692423;
    12'd356: brom_out <= 64'd7165177354826917919;
    12'd357: brom_out <= 64'd4725131077213082099;
    12'd358: brom_out <= 64'd4775626447522085743;
    12'd359: brom_out <= 64'd1916515140755117009;
    12'd360: brom_out <= 64'd6830224072405769937;
    12'd361: brom_out <= 64'd2808578547489358648;
    12'd362: brom_out <= 64'd618886602539794362;
    12'd363: brom_out <= 64'd1761342988433268291;
    12'd364: brom_out <= 64'd7714199699155013517;
    12'd365: brom_out <= 64'd3996172246387663894;
    12'd366: brom_out <= 64'd2407720705974175913;
    12'd367: brom_out <= 64'd845470432081847981;
    12'd368: brom_out <= 64'd5280924731336249208;
    12'd369: brom_out <= 64'd3329477252043532103;
    12'd370: brom_out <= 64'd3865063596590668288;
    12'd371: brom_out <= 64'd896167249461179905;
    12'd372: brom_out <= 64'd6471313754452443304;
    12'd373: brom_out <= 64'd3638579844687192665;
    12'd374: brom_out <= 64'd2648390390780297563;
    12'd375: brom_out <= 64'd4387737789175049378;
    12'd376: brom_out <= 64'd8317572375524300316;
    12'd377: brom_out <= 64'd5053470255903482936;
    12'd378: brom_out <= 64'd9077715168500288810;
    12'd379: brom_out <= 64'd4707096022686776602;
    12'd380: brom_out <= 64'd312660602138865546;
    12'd381: brom_out <= 64'd2837572154281486060;
    12'd382: brom_out <= 64'd2656903131205044847;
    12'd383: brom_out <= 64'd3493841106941144062;
    12'd384: brom_out <= 64'd2744452647294120104;
    12'd385: brom_out <= 64'd5741560898333872640;
    12'd386: brom_out <= 64'd6342775745326442690;
    12'd387: brom_out <= 64'd173655705977138166;
    12'd388: brom_out <= 64'd6767531993306740896;
    12'd389: brom_out <= 64'd510778123162113765;
    12'd390: brom_out <= 64'd6215284701141802918;
    12'd391: brom_out <= 64'd3211346384050301884;
    12'd392: brom_out <= 64'd1742812217555359732;
    12'd393: brom_out <= 64'd6854381567485351737;
    12'd394: brom_out <= 64'd8393653348518333136;
    12'd395: brom_out <= 64'd1414924604129327855;
    12'd396: brom_out <= 64'd3031511680625118659;
    12'd397: brom_out <= 64'd2873657964438583670;
    12'd398: brom_out <= 64'd358825370995750317;
    12'd399: brom_out <= 64'd8388106925642512458;
    12'd400: brom_out <= 64'd4140910720896213055;
    12'd401: brom_out <= 64'd8103768861308718277;
    12'd402: brom_out <= 64'd252340140504241693;
    12'd403: brom_out <= 64'd593580925066186157;
    12'd404: brom_out <= 64'd968670888740781630;
    12'd405: brom_out <= 64'd2825139004329249913;
    12'd406: brom_out <= 64'd7000975899906338725;
    12'd407: brom_out <= 64'd6308865885984590979;
    12'd408: brom_out <= 64'd2311906112180134053;
    12'd409: brom_out <= 64'd4883220479030700178;
    12'd410: brom_out <= 64'd5228929855922500733;
    12'd411: brom_out <= 64'd7570526456457641251;
    12'd412: brom_out <= 64'd5568347348984606631;
    12'd413: brom_out <= 64'd5002301190491438894;
    12'd414: brom_out <= 64'd4330359984991849878;
    12'd415: brom_out <= 64'd278593195830713010;
    12'd416: brom_out <= 64'd3566650897421823420;
    12'd417: brom_out <= 64'd8135274128922892346;
    12'd418: brom_out <= 64'd2706495310779358545;
    12'd419: brom_out <= 64'd6415299222229944443;
    12'd420: brom_out <= 64'd3336750589328840424;
    12'd421: brom_out <= 64'd3716552132217110193;
    12'd422: brom_out <= 64'd7347039844890166366;
    12'd423: brom_out <= 64'd5180232757422409372;
    12'd424: brom_out <= 64'd8733601048999551042;
    12'd425: brom_out <= 64'd8324849038535828029;
    12'd426: brom_out <= 64'd2845549674339093937;
    12'd427: brom_out <= 64'd6996020526618061881;
    12'd428: brom_out <= 64'd729772350383044083;
    12'd429: brom_out <= 64'd3915932020588743220;
    12'd430: brom_out <= 64'd3598529100556018319;
    12'd431: brom_out <= 64'd8533562963389274913;
    12'd432: brom_out <= 64'd6087797337627498753;
    12'd433: brom_out <= 64'd7245595689315409177;
    12'd434: brom_out <= 64'd3654050244854092979;
    12'd435: brom_out <= 64'd8795081828844088731;
    12'd436: brom_out <= 64'd3947696658880618879;
    12'd437: brom_out <= 64'd2780299123311505812;
    12'd438: brom_out <= 64'd7384027011076284535;
    12'd439: brom_out <= 64'd8316279961577302123;
    12'd440: brom_out <= 64'd3434499868985367883;
    12'd441: brom_out <= 64'd3368981121140762329;
    12'd442: brom_out <= 64'd7333818336311565394;
    12'd443: brom_out <= 64'd1750734422805878689;
    12'd444: brom_out <= 64'd8426758779995803383;
    12'd445: brom_out <= 64'd5344604246702031166;
    12'd446: brom_out <= 64'd4017523678350215346;
    12'd447: brom_out <= 64'd2515265228315524440;
    12'd448: brom_out <= 64'd182682343992890333;
    12'd449: brom_out <= 64'd2434563547729207815;
    12'd450: brom_out <= 64'd1883529900336181911;
    12'd451: brom_out <= 64'd2646856009684351864;
    12'd452: brom_out <= 64'd7194983095963719101;
    12'd453: brom_out <= 64'd697957057266428801;
    12'd454: brom_out <= 64'd986365697039853159;
    12'd455: brom_out <= 64'd536607828934758731;
    12'd456: brom_out <= 64'd6675825266329303765;
    12'd457: brom_out <= 64'd9090306241429410261;
    12'd458: brom_out <= 64'd8986601181143710913;
    12'd459: brom_out <= 64'd8089394679902215935;
    12'd460: brom_out <= 64'd8460018361360185973;
    12'd461: brom_out <= 64'd2380034695425169273;
    12'd462: brom_out <= 64'd389354374995615063;
    12'd463: brom_out <= 64'd6566216460598472635;
    12'd464: brom_out <= 64'd468750263104091266;
    12'd465: brom_out <= 64'd2602492081671009787;
    12'd466: brom_out <= 64'd5069373902976902646;
    12'd467: brom_out <= 64'd7927981107379664984;
    12'd468: brom_out <= 64'd5420261389387350880;
    12'd469: brom_out <= 64'd3951152817165964152;
    12'd470: brom_out <= 64'd3017013952813635026;
    12'd471: brom_out <= 64'd3869731669958325174;
    12'd472: brom_out <= 64'd726004773705388864;
    12'd473: brom_out <= 64'd8769091076063025201;
    12'd474: brom_out <= 64'd2610951065952498122;
    12'd475: brom_out <= 64'd7637623102342728356;
    12'd476: brom_out <= 64'd5089878201004960929;
    12'd477: brom_out <= 64'd1569219540301850966;
    12'd478: brom_out <= 64'd7615006295646606520;
    12'd479: brom_out <= 64'd3160635471707226272;
    12'd480: brom_out <= 64'd223404716486023586;
    12'd481: brom_out <= 64'd3706700945489471632;
    12'd482: brom_out <= 64'd1973993570640611291;
    12'd483: brom_out <= 64'd2764856702008527834;
    12'd484: brom_out <= 64'd8235702062124918051;
    12'd485: brom_out <= 64'd6556417574592629401;
    12'd486: brom_out <= 64'd3677374443393723809;
    12'd487: brom_out <= 64'd6822345754583133085;
    12'd488: brom_out <= 64'd2733301067908650870;
    12'd489: brom_out <= 64'd917876077449815305;
    12'd490: brom_out <= 64'd6961232999305020198;
    12'd491: brom_out <= 64'd3440561098919621235;
    12'd492: brom_out <= 64'd1792709974759605982;
    12'd493: brom_out <= 64'd2842470023349595306;
    12'd494: brom_out <= 64'd8019699858674724799;
    12'd495: brom_out <= 64'd7709323644631441076;
    12'd496: brom_out <= 64'd1905920383967759311;
    12'd497: brom_out <= 64'd2780935500684640213;
    12'd498: brom_out <= 64'd5933378338637651478;
    12'd499: brom_out <= 64'd7174739148905575139;
    12'd500: brom_out <= 64'd1752308657048405057;
    12'd501: brom_out <= 64'd3210810410400165574;
    12'd502: brom_out <= 64'd3225264907696276887;
    12'd503: brom_out <= 64'd7344592155860321103;
    12'd504: brom_out <= 64'd693585480357793584;
    12'd505: brom_out <= 64'd5218209040359175169;
    12'd506: brom_out <= 64'd2063677978347548225;
    12'd507: brom_out <= 64'd6115489986575897354;
    12'd508: brom_out <= 64'd7882813018361175933;
    12'd509: brom_out <= 64'd1179590064578720702;
    12'd510: brom_out <= 64'd5061162541301689679;
    12'd511: brom_out <= 64'd5361409663241698187;
    12'd512: brom_out <= 64'd7782386661391366851;
    12'd513: brom_out <= 64'd4861521596590590371;
    12'd514: brom_out <= 64'd8649034445575836908;
    12'd515: brom_out <= 64'd5772687985190368250;
    12'd516: brom_out <= 64'd4381943236453725692;
    12'd517: brom_out <= 64'd3004304654259458127;
    12'd518: brom_out <= 64'd7660778639122281056;
    12'd519: brom_out <= 64'd2835112485135642119;
    12'd520: brom_out <= 64'd2914409323037758834;
    12'd521: brom_out <= 64'd5902160220424771054;
    12'd522: brom_out <= 64'd2585785321548883329;
    12'd523: brom_out <= 64'd1280864215456741565;
    12'd524: brom_out <= 64'd7223163705147076029;
    12'd525: brom_out <= 64'd5481478239653743848;
    12'd526: brom_out <= 64'd8889982071561254404;
    12'd527: brom_out <= 64'd4742566862685097890;
    12'd528: brom_out <= 64'd260052644455523851;
    12'd529: brom_out <= 64'd5559340203372562265;
    12'd530: brom_out <= 64'd6178586593570909300;
    12'd531: brom_out <= 64'd383569141675230395;
    12'd532: brom_out <= 64'd7703760226344578495;
    12'd533: brom_out <= 64'd7508954397386637171;
    12'd534: brom_out <= 64'd2920703367342825301;
    12'd535: brom_out <= 64'd4314847810778816634;
    12'd536: brom_out <= 64'd5652578911009487073;
    12'd537: brom_out <= 64'd9090901240053814193;
    12'd538: brom_out <= 64'd5494996150964866550;
    12'd539: brom_out <= 64'd2118171809324516391;
    12'd540: brom_out <= 64'd3827163200939931713;
    12'd541: brom_out <= 64'd4846498025720647991;
    12'd542: brom_out <= 64'd6510579114601412178;
    12'd543: brom_out <= 64'd7875674622945296174;
    12'd544: brom_out <= 64'd6563344806124755260;
    12'd545: brom_out <= 64'd357276879597893652;
    12'd546: brom_out <= 64'd4124502043139193191;
    12'd547: brom_out <= 64'd6402708749684371457;
    12'd548: brom_out <= 64'd1272215553149008059;
    12'd549: brom_out <= 64'd3539124130597804203;
    12'd550: brom_out <= 64'd4418867056245053493;
    12'd551: brom_out <= 64'd899873894843140087;
    12'd552: brom_out <= 64'd6646628485672871357;
    12'd553: brom_out <= 64'd5885151912454382059;
    12'd554: brom_out <= 64'd6637876692475766041;
    12'd555: brom_out <= 64'd6331760249075063680;
    12'd556: brom_out <= 64'd5208999536819633961;
    12'd557: brom_out <= 64'd4016637484630545084;
    12'd558: brom_out <= 64'd8295305584225460712;
    12'd559: brom_out <= 64'd8277213969632331446;
    12'd560: brom_out <= 64'd6645599729598090252;
    12'd561: brom_out <= 64'd5687432574726921941;
    12'd562: brom_out <= 64'd6624887430223663875;
    12'd563: brom_out <= 64'd8837685408255542790;
    12'd564: brom_out <= 64'd4537650892888119940;
    12'd565: brom_out <= 64'd5346815058652110229;
    12'd566: brom_out <= 64'd4755790540754072763;
    12'd567: brom_out <= 64'd6479702173734099720;
    12'd568: brom_out <= 64'd8138269547828166757;
    12'd569: brom_out <= 64'd570396892100945517;
    12'd570: brom_out <= 64'd1415681576088315011;
    12'd571: brom_out <= 64'd144378385688768922;
    12'd572: brom_out <= 64'd757825782309468411;
    12'd573: brom_out <= 64'd8789340643629732329;
    12'd574: brom_out <= 64'd1762743433048436351;
    12'd575: brom_out <= 64'd3950042927482149122;
    12'd576: brom_out <= 64'd4252522336577894479;
    12'd577: brom_out <= 64'd6633372610416034838;
    12'd578: brom_out <= 64'd266645960251819394;
    12'd579: brom_out <= 64'd5392400538560766981;
    12'd580: brom_out <= 64'd3312612269342758847;
    12'd581: brom_out <= 64'd7630847746185305890;
    12'd582: brom_out <= 64'd2825076588319283267;
    12'd583: brom_out <= 64'd2359484724038118515;
    12'd584: brom_out <= 64'd1703041376499034069;
    12'd585: brom_out <= 64'd7335081421900557064;
    12'd586: brom_out <= 64'd5683902871355065813;
    12'd587: brom_out <= 64'd6487128415723378099;
    12'd588: brom_out <= 64'd6199847152455021322;
    12'd589: brom_out <= 64'd1383247826649431236;
    12'd590: brom_out <= 64'd8104036971331596159;
    12'd591: brom_out <= 64'd7974999663469099555;
    12'd592: brom_out <= 64'd6497957974742993816;
    12'd593: brom_out <= 64'd3776506990065351584;
    12'd594: brom_out <= 64'd8889491850487708094;
    12'd595: brom_out <= 64'd4141239322453315414;
    12'd596: brom_out <= 64'd1821886755871307236;
    12'd597: brom_out <= 64'd8715100417820853311;
    12'd598: brom_out <= 64'd5156989881753429046;
    12'd599: brom_out <= 64'd4482537834370070864;
    12'd600: brom_out <= 64'd5225646594927518733;
    12'd601: brom_out <= 64'd67401699748090272;
    12'd602: brom_out <= 64'd5931022987791557319;
    12'd603: brom_out <= 64'd4699734272960338456;
    12'd604: brom_out <= 64'd6566154634083039334;
    12'd605: brom_out <= 64'd4360439637528448395;
    12'd606: brom_out <= 64'd669990282373323421;
    12'd607: brom_out <= 64'd5467175375755644593;
    12'd608: brom_out <= 64'd2354745007350845777;
    12'd609: brom_out <= 64'd2988079441693257309;
    12'd610: brom_out <= 64'd5198736708809929714;
    12'd611: brom_out <= 64'd3117188644789513996;
    12'd612: brom_out <= 64'd4044154711445931232;
    12'd613: brom_out <= 64'd6885942150999194250;
    12'd614: brom_out <= 64'd2262901270999871265;
    12'd615: brom_out <= 64'd405631466855656892;
    12'd616: brom_out <= 64'd625029411171571798;
    12'd617: brom_out <= 64'd7604631713610068798;
    12'd618: brom_out <= 64'd3130627077031053572;
    12'd619: brom_out <= 64'd7536765662607569693;
    12'd620: brom_out <= 64'd3427924839083361097;
    12'd621: brom_out <= 64'd3310540064712897641;
    12'd622: brom_out <= 64'd3928400720823284202;
    12'd623: brom_out <= 64'd4578784551487833397;
    12'd624: brom_out <= 64'd8061509742389722040;
    12'd625: brom_out <= 64'd6893645876070729278;
    12'd626: brom_out <= 64'd6675720426282350721;
    12'd627: brom_out <= 64'd8656427261785063102;
    12'd628: brom_out <= 64'd5166350325806874424;
    12'd629: brom_out <= 64'd7494705496980488295;
    12'd630: brom_out <= 64'd4549668255283525130;
    12'd631: brom_out <= 64'd1828616697192386803;
    12'd632: brom_out <= 64'd899294709301447584;
    12'd633: brom_out <= 64'd5225422576912013343;
    12'd634: brom_out <= 64'd436640780698173692;
    12'd635: brom_out <= 64'd2776116190172420204;
    12'd636: brom_out <= 64'd8685552408988406375;
    12'd637: brom_out <= 64'd7829622159421577334;
    12'd638: brom_out <= 64'd5585989086796763236;
    12'd639: brom_out <= 64'd7914828735397352007;
    12'd640: brom_out <= 64'd8261458594126653870;
    12'd641: brom_out <= 64'd5739240464631810613;
    12'd642: brom_out <= 64'd4181095021586080784;
    12'd643: brom_out <= 64'd6186822681953179904;
    12'd644: brom_out <= 64'd6107347413120717643;
    12'd645: brom_out <= 64'd6981296114916617638;
    12'd646: brom_out <= 64'd4563281169540611095;
    12'd647: brom_out <= 64'd1526222280158972;
    12'd648: brom_out <= 64'd8033750310262675803;
    12'd649: brom_out <= 64'd3570284798044059338;
    12'd650: brom_out <= 64'd3572599133534823185;
    12'd651: brom_out <= 64'd4456009296275881393;
    12'd652: brom_out <= 64'd6053637598988242858;
    12'd653: brom_out <= 64'd7505420653690884274;
    12'd654: brom_out <= 64'd8347053944178179955;
    12'd655: brom_out <= 64'd6215296105112843792;
    12'd656: brom_out <= 64'd4646018347513530828;
    12'd657: brom_out <= 64'd5811154966774866395;
    12'd658: brom_out <= 64'd7355800531901819327;
    12'd659: brom_out <= 64'd3127006036456972358;
    12'd660: brom_out <= 64'd2824161440388823705;
    12'd661: brom_out <= 64'd4365393897616730227;
    12'd662: brom_out <= 64'd1426929766714741589;
    12'd663: brom_out <= 64'd4944513542595457914;
    12'd664: brom_out <= 64'd3724912625745512029;
    12'd665: brom_out <= 64'd4553170381698880374;
    12'd666: brom_out <= 64'd7040172441218270691;
    12'd667: brom_out <= 64'd2678802622163617608;
    12'd668: brom_out <= 64'd680992054214511747;
    12'd669: brom_out <= 64'd5234674833021145037;
    12'd670: brom_out <= 64'd6069141774778254976;
    12'd671: brom_out <= 64'd1599192383156885901;
    12'd672: brom_out <= 64'd3112085083619698235;
    12'd673: brom_out <= 64'd8808466971874321347;
    12'd674: brom_out <= 64'd1742075655550483472;
    12'd675: brom_out <= 64'd1560624357375366680;
    12'd676: brom_out <= 64'd931917372433455172;
    12'd677: brom_out <= 64'd3948779935617512385;
    12'd678: brom_out <= 64'd8513457866454952299;
    12'd679: brom_out <= 64'd8071993320658122545;
    12'd680: brom_out <= 64'd6838354098954707793;
    12'd681: brom_out <= 64'd6452037462833976715;
    12'd682: brom_out <= 64'd3940981814208109053;
    12'd683: brom_out <= 64'd7921735501324498558;
    12'd684: brom_out <= 64'd3017522447692063281;
    12'd685: brom_out <= 64'd1576647487118034598;
    12'd686: brom_out <= 64'd2738988075928486416;
    12'd687: brom_out <= 64'd7328417818605634705;
    12'd688: brom_out <= 64'd7060407982316328557;
    12'd689: brom_out <= 64'd7380059655556803829;
    12'd690: brom_out <= 64'd6537574420544680745;
    12'd691: brom_out <= 64'd7985284825629649381;
    12'd692: brom_out <= 64'd7068134865767266017;
    12'd693: brom_out <= 64'd4384544437249056579;
    12'd694: brom_out <= 64'd5029278047678630553;
    12'd695: brom_out <= 64'd2442215543049826913;
    12'd696: brom_out <= 64'd8061035613661260463;
    12'd697: brom_out <= 64'd1769305370968412801;
    12'd698: brom_out <= 64'd1818887195464307806;
    12'd699: brom_out <= 64'd3668231896105362147;
    12'd700: brom_out <= 64'd1596191628058893204;
    12'd701: brom_out <= 64'd3852766516875788633;
    12'd702: brom_out <= 64'd5476941396846307088;
    12'd703: brom_out <= 64'd1058480063031661059;
    12'd704: brom_out <= 64'd95281317708976622;
    12'd705: brom_out <= 64'd4011203195838380948;
    12'd706: brom_out <= 64'd27725867473174067;
    12'd707: brom_out <= 64'd944892544399607082;
    12'd708: brom_out <= 64'd5767241774841291582;
    12'd709: brom_out <= 64'd7146643211714477250;
    12'd710: brom_out <= 64'd8234010378906857987;
    12'd711: brom_out <= 64'd8738310441896228275;
    12'd712: brom_out <= 64'd437504944868661480;
    12'd713: brom_out <= 64'd1345594068393668289;
    12'd714: brom_out <= 64'd7790278521481987032;
    12'd715: brom_out <= 64'd11091872513553694;
    12'd716: brom_out <= 64'd2458237992137544474;
    12'd717: brom_out <= 64'd7480666283181908954;
    12'd718: brom_out <= 64'd8096484272479559454;
    12'd719: brom_out <= 64'd7045313376099365566;
    12'd720: brom_out <= 64'd3594081468019201941;
    12'd721: brom_out <= 64'd2574614894679130082;
    12'd722: brom_out <= 64'd5412263672042607496;
    12'd723: brom_out <= 64'd952462368163070319;
    12'd724: brom_out <= 64'd8686991881157190307;
    12'd725: brom_out <= 64'd1985359551968673528;
    12'd726: brom_out <= 64'd4675753835282043687;
    12'd727: brom_out <= 64'd7276908357077529473;
    12'd728: brom_out <= 64'd5272909420026529286;
    12'd729: brom_out <= 64'd7041957683143414597;
    12'd730: brom_out <= 64'd7923353732097988637;
    12'd731: brom_out <= 64'd7622846587038404776;
    12'd732: brom_out <= 64'd5866323178725112845;
    12'd733: brom_out <= 64'd5200255370324995803;
    12'd734: brom_out <= 64'd4967626057439603150;
    12'd735: brom_out <= 64'd4409427483205928698;
    12'd736: brom_out <= 64'd7504794892223181970;
    12'd737: brom_out <= 64'd7112929143432610457;
    12'd738: brom_out <= 64'd6857070551449887647;
    12'd739: brom_out <= 64'd6550567352823378811;
    12'd740: brom_out <= 64'd7990782566459026937;
    12'd741: brom_out <= 64'd3512327954730964416;
    12'd742: brom_out <= 64'd2756726733978479127;
    12'd743: brom_out <= 64'd6627709141254412355;
    12'd744: brom_out <= 64'd1207092097272907855;
    12'd745: brom_out <= 64'd8714591519982473863;
    12'd746: brom_out <= 64'd2202922525939669635;
    12'd747: brom_out <= 64'd1742247754033219684;
    12'd748: brom_out <= 64'd4267532708699862748;
    12'd749: brom_out <= 64'd6325751102943649754;
    12'd750: brom_out <= 64'd9126508312536893339;
    12'd751: brom_out <= 64'd7276369704671830683;
    12'd752: brom_out <= 64'd3936456730853119832;
    12'd753: brom_out <= 64'd6316914292526049085;
    12'd754: brom_out <= 64'd671388122160422741;
    12'd755: brom_out <= 64'd7721993641687260771;
    12'd756: brom_out <= 64'd6593077827335687009;
    12'd757: brom_out <= 64'd1471472388324251922;
    12'd758: brom_out <= 64'd4840954178999118923;
    12'd759: brom_out <= 64'd3206943792237108235;
    12'd760: brom_out <= 64'd3869156205775182321;
    12'd761: brom_out <= 64'd3079940288112575077;
    12'd762: brom_out <= 64'd6846128385768296431;
    12'd763: brom_out <= 64'd26364125632882708;
    12'd764: brom_out <= 64'd2919108040339750211;
    12'd765: brom_out <= 64'd8768781517050275053;
    12'd766: brom_out <= 64'd6955996116910048576;
    12'd767: brom_out <= 64'd2459613877402660323;
    12'd768: brom_out <= 64'd3666700039899848147;
    12'd769: brom_out <= 64'd6902448893183730201;
    12'd770: brom_out <= 64'd2624606603770530868;
    12'd771: brom_out <= 64'd6670734812323184165;
    12'd772: brom_out <= 64'd7280238195358008995;
    12'd773: brom_out <= 64'd2015983383132894781;
    12'd774: brom_out <= 64'd2466974359874510230;
    12'd775: brom_out <= 64'd6460324180094717038;
    12'd776: brom_out <= 64'd6844075998943291247;
    12'd777: brom_out <= 64'd6033708933034981867;
    12'd778: brom_out <= 64'd9112820884944911520;
    12'd779: brom_out <= 64'd9122891899647476238;
    12'd780: brom_out <= 64'd4827416146413489003;
    12'd781: brom_out <= 64'd1525777051077072050;
    12'd782: brom_out <= 64'd8336562908643181499;
    12'd783: brom_out <= 64'd6685683477184525655;
    12'd784: brom_out <= 64'd6165347185232428134;
    12'd785: brom_out <= 64'd319725465409657507;
    12'd786: brom_out <= 64'd2527881211643169611;
    12'd787: brom_out <= 64'd2035157007536029201;
    12'd788: brom_out <= 64'd5444954182365675077;
    12'd789: brom_out <= 64'd2856848174308624223;
    12'd790: brom_out <= 64'd4210509491007543576;
    12'd791: brom_out <= 64'd3985754481246278600;
    12'd792: brom_out <= 64'd1207978512304215843;
    12'd793: brom_out <= 64'd6426530318111945989;
    12'd794: brom_out <= 64'd6839147203842741647;
    12'd795: brom_out <= 64'd1099540133965673030;
    12'd796: brom_out <= 64'd8370814366380482311;
    12'd797: brom_out <= 64'd9175914659917467912;
    12'd798: brom_out <= 64'd5821644811909952191;
    12'd799: brom_out <= 64'd2878034258543693224;
    12'd800: brom_out <= 64'd4238249638059871551;
    12'd801: brom_out <= 64'd7708655880151707474;
    12'd802: brom_out <= 64'd2695807627030083465;
    12'd803: brom_out <= 64'd1346451435635629720;
    12'd804: brom_out <= 64'd7390346186579725385;
    12'd805: brom_out <= 64'd9089560507989965207;
    12'd806: brom_out <= 64'd8267751919188170351;
    12'd807: brom_out <= 64'd6213190605695911440;
    12'd808: brom_out <= 64'd6507088774975524892;
    12'd809: brom_out <= 64'd4410029091311437334;
    12'd810: brom_out <= 64'd6359903742957886409;
    12'd811: brom_out <= 64'd4654745623883232599;
    12'd812: brom_out <= 64'd2197487004130961575;
    12'd813: brom_out <= 64'd2829576829854501102;
    12'd814: brom_out <= 64'd8940771018146404979;
    12'd815: brom_out <= 64'd4354317671001826892;
    12'd816: brom_out <= 64'd4561515202707775996;
    12'd817: brom_out <= 64'd432118055352980039;
    12'd818: brom_out <= 64'd6089338024589188016;
    12'd819: brom_out <= 64'd7565980322032079733;
    12'd820: brom_out <= 64'd5621318752886328;
    12'd821: brom_out <= 64'd2081185830936091222;
    12'd822: brom_out <= 64'd6700248938855750088;
    12'd823: brom_out <= 64'd6109644353229462220;
    12'd824: brom_out <= 64'd4127725377931775362;
    12'd825: brom_out <= 64'd3445536536338924127;
    12'd826: brom_out <= 64'd8039663376801308076;
    12'd827: brom_out <= 64'd2039924189795129333;
    12'd828: brom_out <= 64'd1762152160220190022;
    12'd829: brom_out <= 64'd6227684377220662635;
    12'd830: brom_out <= 64'd3460699204374494731;
    12'd831: brom_out <= 64'd2507386577908709969;
    12'd832: brom_out <= 64'd9171435364368087656;
    12'd833: brom_out <= 64'd2704736918382890252;
    12'd834: brom_out <= 64'd6867932455866769948;
    12'd835: brom_out <= 64'd4733223220944963107;
    12'd836: brom_out <= 64'd89191171625464338;
    12'd837: brom_out <= 64'd2996845867260708288;
    12'd838: brom_out <= 64'd1330423127781123172;
    12'd839: brom_out <= 64'd8813447416130232538;
    12'd840: brom_out <= 64'd3041920256613138472;
    12'd841: brom_out <= 64'd5287685692033182571;
    12'd842: brom_out <= 64'd1554685205797863112;
    12'd843: brom_out <= 64'd2679623975545059377;
    12'd844: brom_out <= 64'd8619418134468106589;
    12'd845: brom_out <= 64'd866252214217421753;
    12'd846: brom_out <= 64'd3744644079555530802;
    12'd847: brom_out <= 64'd4835801822145010876;
    12'd848: brom_out <= 64'd8634953690816838135;
    12'd849: brom_out <= 64'd4649853355221802222;
    12'd850: brom_out <= 64'd981653074263351650;
    12'd851: brom_out <= 64'd5821311771166244451;
    12'd852: brom_out <= 64'd5607126821066373889;
    12'd853: brom_out <= 64'd1556875117719560478;
    12'd854: brom_out <= 64'd5227909491507430272;
    12'd855: brom_out <= 64'd7808349424018495852;
    12'd856: brom_out <= 64'd4636341520660054868;
    12'd857: brom_out <= 64'd8961140586297088736;
    12'd858: brom_out <= 64'd6807079627032911582;
    12'd859: brom_out <= 64'd7084188348831055435;
    12'd860: brom_out <= 64'd5031374273336242327;
    12'd861: brom_out <= 64'd375186616369405533;
    12'd862: brom_out <= 64'd610804669399733493;
    12'd863: brom_out <= 64'd3025306996498679989;
    12'd864: brom_out <= 64'd6737329518480497135;
    12'd865: brom_out <= 64'd2048220758058706870;
    12'd866: brom_out <= 64'd3189897571657284634;
    12'd867: brom_out <= 64'd768889390292241765;
    12'd868: brom_out <= 64'd2647786732026981346;
    12'd869: brom_out <= 64'd36752078914957114;
    12'd870: brom_out <= 64'd247805208039003867;
    12'd871: brom_out <= 64'd2511839478159507331;
    12'd872: brom_out <= 64'd2516463966353163527;
    12'd873: brom_out <= 64'd4205791328057774404;
    12'd874: brom_out <= 64'd1979255590725765209;
    12'd875: brom_out <= 64'd1179978746940840805;
    12'd876: brom_out <= 64'd1648540804641590701;
    12'd877: brom_out <= 64'd9000560894531380343;
    12'd878: brom_out <= 64'd799001452467389122;
    12'd879: brom_out <= 64'd6077440687542564946;
    12'd880: brom_out <= 64'd1366069914788878450;
    12'd881: brom_out <= 64'd8488803381524692255;
    12'd882: brom_out <= 64'd2304688208552581358;
    12'd883: brom_out <= 64'd3782017943009885866;
    12'd884: brom_out <= 64'd5881118486570837651;
    12'd885: brom_out <= 64'd4427602785075522478;
    12'd886: brom_out <= 64'd152427030840984604;
    12'd887: brom_out <= 64'd5078921445156716018;
    12'd888: brom_out <= 64'd9083664109308128459;
    12'd889: brom_out <= 64'd1845931253922829248;
    12'd890: brom_out <= 64'd3306135986659390567;
    12'd891: brom_out <= 64'd2925974740967275136;
    12'd892: brom_out <= 64'd8105079806250145642;
    12'd893: brom_out <= 64'd2988226832345877022;
    12'd894: brom_out <= 64'd1435161344878474098;
    12'd895: brom_out <= 64'd8457738163840186981;
    12'd896: brom_out <= 64'd4402385349865443935;
    12'd897: brom_out <= 64'd8226036132022963627;
    12'd898: brom_out <= 64'd4255379659518795183;
    12'd899: brom_out <= 64'd6411389752420834287;
    12'd900: brom_out <= 64'd3601109703153377607;
    12'd901: brom_out <= 64'd2609445345925526117;
    12'd902: brom_out <= 64'd5393687233907933846;
    12'd903: brom_out <= 64'd4231299252631786363;
    12'd904: brom_out <= 64'd7611455445751931128;
    12'd905: brom_out <= 64'd5556737181015255713;
    12'd906: brom_out <= 64'd3178783619418943918;
    12'd907: brom_out <= 64'd6666399481015416211;
    12'd908: brom_out <= 64'd1476606023428051712;
    12'd909: brom_out <= 64'd4897891012526249384;
    12'd910: brom_out <= 64'd807621101160052175;
    12'd911: brom_out <= 64'd4485097006786027744;
    12'd912: brom_out <= 64'd3961328919819112353;
    12'd913: brom_out <= 64'd7270855825469751732;
    12'd914: brom_out <= 64'd1870792994676811958;
    12'd915: brom_out <= 64'd4178561717271544320;
    12'd916: brom_out <= 64'd5330596359306770007;
    12'd917: brom_out <= 64'd4994830263320322381;
    12'd918: brom_out <= 64'd3888759199275104826;
    12'd919: brom_out <= 64'd6358460373818083425;
    12'd920: brom_out <= 64'd7793709421929414301;
    12'd921: brom_out <= 64'd7066411863153210917;
    12'd922: brom_out <= 64'd8239775268200818068;
    12'd923: brom_out <= 64'd2577794354245569325;
    12'd924: brom_out <= 64'd7364279298402482039;
    12'd925: brom_out <= 64'd4990831297253965132;
    12'd926: brom_out <= 64'd7187784025358661201;
    12'd927: brom_out <= 64'd8837090426427861905;
    12'd928: brom_out <= 64'd7892893190033330700;
    12'd929: brom_out <= 64'd5837236979066677584;
    12'd930: brom_out <= 64'd3209619641628172834;
    12'd931: brom_out <= 64'd7633757610897567398;
    12'd932: brom_out <= 64'd201270148177865980;
    12'd933: brom_out <= 64'd2812886942652402345;
    12'd934: brom_out <= 64'd2132564876249104045;
    12'd935: brom_out <= 64'd829786685533664686;
    12'd936: brom_out <= 64'd4158304906226181360;
    12'd937: brom_out <= 64'd8339234857201480490;
    12'd938: brom_out <= 64'd8109255189159764048;
    12'd939: brom_out <= 64'd2037752842496234735;
    12'd940: brom_out <= 64'd6565289806182052066;
    12'd941: brom_out <= 64'd4793923028636351289;
    12'd942: brom_out <= 64'd5786909569893455239;
    12'd943: brom_out <= 64'd1246867284200325980;
    12'd944: brom_out <= 64'd8875392094220290763;
    12'd945: brom_out <= 64'd8459532325918774522;
    12'd946: brom_out <= 64'd560707250059269947;
    12'd947: brom_out <= 64'd6481694119177686866;
    12'd948: brom_out <= 64'd4119638043528018860;
    12'd949: brom_out <= 64'd6206251482753171757;
    12'd950: brom_out <= 64'd8870261372249595655;
    12'd951: brom_out <= 64'd6165341452860093577;
    12'd952: brom_out <= 64'd8524663551246023401;
    12'd953: brom_out <= 64'd1614715635848808903;
    12'd954: brom_out <= 64'd267001868020741669;
    12'd955: brom_out <= 64'd5881703684718594878;
    12'd956: brom_out <= 64'd2992569522693031963;
    12'd957: brom_out <= 64'd6805038745224127631;
    12'd958: brom_out <= 64'd4818694961486043108;
    12'd959: brom_out <= 64'd5860526560614714467;
    12'd960: brom_out <= 64'd1301058986836242658;
    12'd961: brom_out <= 64'd2046057320205376781;
    12'd962: brom_out <= 64'd7288514495394200147;
    12'd963: brom_out <= 64'd2633859063286017972;
    12'd964: brom_out <= 64'd9008652145339594081;
    12'd965: brom_out <= 64'd8458397413255347953;
    12'd966: brom_out <= 64'd9003992428561474784;
    12'd967: brom_out <= 64'd6396892344171279300;
    12'd968: brom_out <= 64'd8467731552125190747;
    12'd969: brom_out <= 64'd3577344067180045365;
    12'd970: brom_out <= 64'd9060560875587670594;
    12'd971: brom_out <= 64'd3801514624142414422;
    12'd972: brom_out <= 64'd4382892675974943446;
    12'd973: brom_out <= 64'd4149902099744216290;
    12'd974: brom_out <= 64'd7066430919226304905;
    12'd975: brom_out <= 64'd6334509964978317045;
    12'd976: brom_out <= 64'd6889211782122528516;
    12'd977: brom_out <= 64'd2150239118104650937;
    12'd978: brom_out <= 64'd5746120609323938049;
    12'd979: brom_out <= 64'd6541337151798288460;
    12'd980: brom_out <= 64'd3084270353954939594;
    12'd981: brom_out <= 64'd4319368292303648262;
    12'd982: brom_out <= 64'd427711520458827573;
    12'd983: brom_out <= 64'd8844779975228976583;
    12'd984: brom_out <= 64'd235928975280521441;
    12'd985: brom_out <= 64'd2613405612301128147;
    12'd986: brom_out <= 64'd4154410606352405184;
    12'd987: brom_out <= 64'd9068096702955046917;
    12'd988: brom_out <= 64'd4178188816799367836;
    12'd989: brom_out <= 64'd2142244415983486190;
    12'd990: brom_out <= 64'd8979329132321310905;
    12'd991: brom_out <= 64'd6967090839982818812;
    12'd992: brom_out <= 64'd4190939924922756337;
    12'd993: brom_out <= 64'd5676361374244060971;
    12'd994: brom_out <= 64'd9033577227275030048;
    12'd995: brom_out <= 64'd8450886564708926769;
    12'd996: brom_out <= 64'd2689097136219244759;
    12'd997: brom_out <= 64'd3600413203762509257;
    12'd998: brom_out <= 64'd3948633174989000328;
    12'd999: brom_out <= 64'd3755891007880143387;
    12'd1000: brom_out <= 64'd1776169442401324753;
    12'd1001: brom_out <= 64'd4405927027337897707;
    12'd1002: brom_out <= 64'd359322144804628539;
    12'd1003: brom_out <= 64'd6698642343086080125;
    12'd1004: brom_out <= 64'd5145517706759223898;
    12'd1005: brom_out <= 64'd1662890316899717972;
    12'd1006: brom_out <= 64'd5380475214395068961;
    12'd1007: brom_out <= 64'd6674765443416448252;
    12'd1008: brom_out <= 64'd1079581639635537229;
    12'd1009: brom_out <= 64'd3257049769028043096;
    12'd1010: brom_out <= 64'd1975844918861245996;
    12'd1011: brom_out <= 64'd2753051010196344335;
    12'd1012: brom_out <= 64'd5589004524259874951;
    12'd1013: brom_out <= 64'd7686967573819799816;
    12'd1014: brom_out <= 64'd8837279335233063974;
    12'd1015: brom_out <= 64'd8479001584131948299;
    12'd1016: brom_out <= 64'd4009441159250921872;
    12'd1017: brom_out <= 64'd4942129846177841682;
    12'd1018: brom_out <= 64'd6181169933655709384;
    12'd1019: brom_out <= 64'd2088737596298706012;
    12'd1020: brom_out <= 64'd1187360867394053595;
    12'd1021: brom_out <= 64'd3169187917214977042;
    12'd1022: brom_out <= 64'd4094156051496113580;
    12'd1023: brom_out <= 64'd5812672108857599105;
    12'd1024: brom_out <= 64'd3524599538144401835;
    12'd1025: brom_out <= 64'd965865660521274904;
    12'd1026: brom_out <= 64'd6038219084579328985;
    12'd1027: brom_out <= 64'd4592595758117140191;
    12'd1028: brom_out <= 64'd8825067894575323629;
    12'd1029: brom_out <= 64'd3346724334594068778;
    12'd1030: brom_out <= 64'd5196642866436430279;
    12'd1031: brom_out <= 64'd7267243829075110462;
    12'd1032: brom_out <= 64'd4243922567581545872;
    12'd1033: brom_out <= 64'd4962202444033985523;
    12'd1034: brom_out <= 64'd3678639522642170811;
    12'd1035: brom_out <= 64'd4699341332070757189;
    12'd1036: brom_out <= 64'd884291909185288083;
    12'd1037: brom_out <= 64'd7195166790530456084;
    12'd1038: brom_out <= 64'd7128421414828377760;
    12'd1039: brom_out <= 64'd4036162231626469298;
    12'd1040: brom_out <= 64'd1312032635293907300;
    12'd1041: brom_out <= 64'd4014799508541499699;
    12'd1042: brom_out <= 64'd7558797298569106217;
    12'd1043: brom_out <= 64'd2236080304131579697;
    12'd1044: brom_out <= 64'd2208983202347601940;
    12'd1045: brom_out <= 64'd8893574271825646043;
    12'd1046: brom_out <= 64'd1845434832961287151;
    12'd1047: brom_out <= 64'd933077087322545712;
    12'd1048: brom_out <= 64'd4883309178694173302;
    12'd1049: brom_out <= 64'd5704817086217644123;
    12'd1050: brom_out <= 64'd5204926216551210872;
    12'd1051: brom_out <= 64'd6200385498913318034;
    12'd1052: brom_out <= 64'd7082252839057205732;
    12'd1053: brom_out <= 64'd210419244933660052;
    12'd1054: brom_out <= 64'd6503085852836274346;
    12'd1055: brom_out <= 64'd1544824365766875241;
    12'd1056: brom_out <= 64'd941177897218823962;
    12'd1057: brom_out <= 64'd7389367459254262663;
    12'd1058: brom_out <= 64'd5365720439767022829;
    12'd1059: brom_out <= 64'd2255462934494463142;
    12'd1060: brom_out <= 64'd4536966134794454621;
    12'd1061: brom_out <= 64'd1385947144974908023;
    12'd1062: brom_out <= 64'd619338145319270643;
    12'd1063: brom_out <= 64'd6791000566943613855;
    12'd1064: brom_out <= 64'd823754380868015806;
    12'd1065: brom_out <= 64'd5709651044590000246;
    12'd1066: brom_out <= 64'd804601355462899423;
    12'd1067: brom_out <= 64'd7082077200405620635;
    12'd1068: brom_out <= 64'd8905793174997083851;
    12'd1069: brom_out <= 64'd635036423699835615;
    12'd1070: brom_out <= 64'd7076613822757551988;
    12'd1071: brom_out <= 64'd753458034391468420;
    12'd1072: brom_out <= 64'd7896337347699643758;
    12'd1073: brom_out <= 64'd366757094310288330;
    12'd1074: brom_out <= 64'd2050583595339069286;
    12'd1075: brom_out <= 64'd4083343559744628073;
    12'd1076: brom_out <= 64'd7275280601212547141;
    12'd1077: brom_out <= 64'd6276005299585931277;
    12'd1078: brom_out <= 64'd5848149142182723081;
    12'd1079: brom_out <= 64'd7405531063152648609;
    12'd1080: brom_out <= 64'd2247898014124480324;
    12'd1081: brom_out <= 64'd2531633857331206109;
    12'd1082: brom_out <= 64'd1951441445411639130;
    12'd1083: brom_out <= 64'd6608021666455320110;
    12'd1084: brom_out <= 64'd4315824744591934752;
    12'd1085: brom_out <= 64'd7384227251435011657;
    12'd1086: brom_out <= 64'd5364611743911052676;
    12'd1087: brom_out <= 64'd3104797388995996590;
    12'd1088: brom_out <= 64'd6855776959140026846;
    12'd1089: brom_out <= 64'd3008739132914375284;
    12'd1090: brom_out <= 64'd1800152208982219194;
    12'd1091: brom_out <= 64'd4536620460504430233;
    12'd1092: brom_out <= 64'd1072795248158240320;
    12'd1093: brom_out <= 64'd3651471097977905112;
    12'd1094: brom_out <= 64'd5592076851950722483;
    12'd1095: brom_out <= 64'd91888639829313925;
    12'd1096: brom_out <= 64'd6092339191021377621;
    12'd1097: brom_out <= 64'd4201276373534048168;
    12'd1098: brom_out <= 64'd6899783450675602801;
    12'd1099: brom_out <= 64'd4354852178817980642;
    12'd1100: brom_out <= 64'd8078584416777687580;
    12'd1101: brom_out <= 64'd8988613599268288848;
    12'd1102: brom_out <= 64'd1396460064938311569;
    12'd1103: brom_out <= 64'd4808499690770491665;
    12'd1104: brom_out <= 64'd770547429306764387;
    12'd1105: brom_out <= 64'd7452564609534301780;
    12'd1106: brom_out <= 64'd8913398684432203431;
    12'd1107: brom_out <= 64'd1589588185396114735;
    12'd1108: brom_out <= 64'd7931311122728956933;
    12'd1109: brom_out <= 64'd4506266599100625746;
    12'd1110: brom_out <= 64'd812033014687402642;
    12'd1111: brom_out <= 64'd3891046209747111995;
    12'd1112: brom_out <= 64'd7775530046837291397;
    12'd1113: brom_out <= 64'd7954176500850726075;
    12'd1114: brom_out <= 64'd6773413460164400989;
    12'd1115: brom_out <= 64'd3544126875777306127;
    12'd1116: brom_out <= 64'd1561735603309602318;
    12'd1117: brom_out <= 64'd564287763593718972;
    12'd1118: brom_out <= 64'd1319625945528114437;
    12'd1119: brom_out <= 64'd653641936569555104;
    12'd1120: brom_out <= 64'd1654143360053197228;
    12'd1121: brom_out <= 64'd6100972164166701452;
    12'd1122: brom_out <= 64'd7009740899173647904;
    12'd1123: brom_out <= 64'd391244183956117656;
    12'd1124: brom_out <= 64'd6658501207946687856;
    12'd1125: brom_out <= 64'd4837928164813805094;
    12'd1126: brom_out <= 64'd1246869919003470948;
    12'd1127: brom_out <= 64'd4556396931413170565;
    12'd1128: brom_out <= 64'd2901067591160354491;
    12'd1129: brom_out <= 64'd7237123114547387231;
    12'd1130: brom_out <= 64'd6956094196580450535;
    12'd1131: brom_out <= 64'd8078096999426657769;
    12'd1132: brom_out <= 64'd6996719195351172105;
    12'd1133: brom_out <= 64'd3042494614533923543;
    12'd1134: brom_out <= 64'd12532349657011920;
    12'd1135: brom_out <= 64'd6323756161825652617;
    12'd1136: brom_out <= 64'd7340614074242873515;
    12'd1137: brom_out <= 64'd419344938408565205;
    12'd1138: brom_out <= 64'd2499939223131857379;
    12'd1139: brom_out <= 64'd8769856015462760900;
    12'd1140: brom_out <= 64'd4405462643572670401;
    12'd1141: brom_out <= 64'd2600721565327225693;
    12'd1142: brom_out <= 64'd3554411748700026067;
    12'd1143: brom_out <= 64'd5105121559920632872;
    12'd1144: brom_out <= 64'd5044677667335809588;
    12'd1145: brom_out <= 64'd855019649065814602;
    12'd1146: brom_out <= 64'd2116795489411995706;
    12'd1147: brom_out <= 64'd8450532263755236763;
    12'd1148: brom_out <= 64'd6192001440112219942;
    12'd1149: brom_out <= 64'd3925032875092237225;
    12'd1150: brom_out <= 64'd4827353238050434248;
    12'd1151: brom_out <= 64'd845949387679313112;
    12'd1152: brom_out <= 64'd1037226495264959765;
    12'd1153: brom_out <= 64'd3184802302563900160;
    12'd1154: brom_out <= 64'd6092418754942118738;
    12'd1155: brom_out <= 64'd1498043933519780510;
    12'd1156: brom_out <= 64'd1304184122061830153;
    12'd1157: brom_out <= 64'd4861844953477305444;
    12'd1158: brom_out <= 64'd5076072023075556729;
    12'd1159: brom_out <= 64'd8385145770674892915;
    12'd1160: brom_out <= 64'd2546715249149327980;
    12'd1161: brom_out <= 64'd1031728823264968702;
    12'd1162: brom_out <= 64'd9077463387344432871;
    12'd1163: brom_out <= 64'd7700144060295659713;
    12'd1164: brom_out <= 64'd5247116371508764185;
    12'd1165: brom_out <= 64'd3582103710376572665;
    12'd1166: brom_out <= 64'd3208657701039362660;
    12'd1167: brom_out <= 64'd4968325785424395217;
    12'd1168: brom_out <= 64'd1945060455200500649;
    12'd1169: brom_out <= 64'd7647775544549925544;
    12'd1170: brom_out <= 64'd4632934557344117998;
    12'd1171: brom_out <= 64'd4249755460971679640;
    12'd1172: brom_out <= 64'd6307520490536919089;
    12'd1173: brom_out <= 64'd6145327616371340629;
    12'd1174: brom_out <= 64'd5656979822188425455;
    12'd1175: brom_out <= 64'd7171380709763832871;
    12'd1176: brom_out <= 64'd3980571863301283620;
    12'd1177: brom_out <= 64'd2895327248236271286;
    12'd1178: brom_out <= 64'd7025921624635260245;
    12'd1179: brom_out <= 64'd7559606478731311905;
    12'd1180: brom_out <= 64'd1279915414899990542;
    12'd1181: brom_out <= 64'd4166692459634219505;
    12'd1182: brom_out <= 64'd282350079186146223;
    12'd1183: brom_out <= 64'd8785704162863890026;
    12'd1184: brom_out <= 64'd2519409300647451668;
    12'd1185: brom_out <= 64'd4488325412383412473;
    12'd1186: brom_out <= 64'd6937670974143645308;
    12'd1187: brom_out <= 64'd6399717363275658235;
    12'd1188: brom_out <= 64'd3434456093458602952;
    12'd1189: brom_out <= 64'd280046794241272709;
    12'd1190: brom_out <= 64'd2925582264698277317;
    12'd1191: brom_out <= 64'd1532519841461757190;
    12'd1192: brom_out <= 64'd8980860614517287927;
    12'd1193: brom_out <= 64'd7353004483382456242;
    12'd1194: brom_out <= 64'd8856043797460319807;
    12'd1195: brom_out <= 64'd6826497808383185357;
    12'd1196: brom_out <= 64'd8942821574826056080;
    12'd1197: brom_out <= 64'd4060323279366876069;
    12'd1198: brom_out <= 64'd1573727348570003143;
    12'd1199: brom_out <= 64'd3461538383816916234;
    12'd1200: brom_out <= 64'd5525258807420722821;
    12'd1201: brom_out <= 64'd568649861241646821;
    12'd1202: brom_out <= 64'd1363262778621793103;
    12'd1203: brom_out <= 64'd4742697653959067366;
    12'd1204: brom_out <= 64'd4484144502716956109;
    12'd1205: brom_out <= 64'd3469576714098428976;
    12'd1206: brom_out <= 64'd1967907399506487696;
    12'd1207: brom_out <= 64'd6906947201749861657;
    12'd1208: brom_out <= 64'd2382835902027319685;
    12'd1209: brom_out <= 64'd7261099267870562601;
    12'd1210: brom_out <= 64'd7830596987955495764;
    12'd1211: brom_out <= 64'd9184156761960620759;
    12'd1212: brom_out <= 64'd3073145352091067037;
    12'd1213: brom_out <= 64'd7172546964820155978;
    12'd1214: brom_out <= 64'd2189336162637014780;
    12'd1215: brom_out <= 64'd4607562414967830263;
    12'd1216: brom_out <= 64'd143040478232822066;
    12'd1217: brom_out <= 64'd1485252593272270883;
    12'd1218: brom_out <= 64'd4267852789840945245;
    12'd1219: brom_out <= 64'd6707927437333985301;
    12'd1220: brom_out <= 64'd9061361895215172237;
    12'd1221: brom_out <= 64'd468324080733551514;
    12'd1222: brom_out <= 64'd4918085894909184471;
    12'd1223: brom_out <= 64'd4598611642296756705;
    12'd1224: brom_out <= 64'd7433084580286989857;
    12'd1225: brom_out <= 64'd5866700892828110188;
    12'd1226: brom_out <= 64'd2389457907874897124;
    12'd1227: brom_out <= 64'd2910226872121544553;
    12'd1228: brom_out <= 64'd9077092935487857308;
    12'd1229: brom_out <= 64'd4799307411913717518;
    12'd1230: brom_out <= 64'd3203935204274517324;
    12'd1231: brom_out <= 64'd38850968059739164;
    12'd1232: brom_out <= 64'd4624281104272904919;
    12'd1233: brom_out <= 64'd2456615652581159166;
    12'd1234: brom_out <= 64'd213881384110140280;
    12'd1235: brom_out <= 64'd9164877232180664454;
    12'd1236: brom_out <= 64'd9032974342355614921;
    12'd1237: brom_out <= 64'd4863773591867402437;
    12'd1238: brom_out <= 64'd5820943596997641184;
    12'd1239: brom_out <= 64'd2336160345686382031;
    12'd1240: brom_out <= 64'd805362609902649459;
    12'd1241: brom_out <= 64'd7633242113754359003;
    12'd1242: brom_out <= 64'd3591956466773264267;
    12'd1243: brom_out <= 64'd3436169704694582004;
    12'd1244: brom_out <= 64'd179191309904241533;
    12'd1245: brom_out <= 64'd9151570473005599210;
    12'd1246: brom_out <= 64'd8967626807078366641;
    12'd1247: brom_out <= 64'd3218248454179245766;
    12'd1248: brom_out <= 64'd531312113401045055;
    12'd1249: brom_out <= 64'd7411062221110083731;
    12'd1250: brom_out <= 64'd7053149561235473502;
    12'd1251: brom_out <= 64'd6714704800367854718;
    12'd1252: brom_out <= 64'd321539602964568364;
    12'd1253: brom_out <= 64'd6044797564155680637;
    12'd1254: brom_out <= 64'd1875475665087908322;
    12'd1255: brom_out <= 64'd600741020216472508;
    12'd1256: brom_out <= 64'd8706280792139117950;
    12'd1257: brom_out <= 64'd6586920412784111395;
    12'd1258: brom_out <= 64'd4352875976613107716;
    12'd1259: brom_out <= 64'd2062454173864398730;
    12'd1260: brom_out <= 64'd1264319546698281601;
    12'd1261: brom_out <= 64'd7043989661891023753;
    12'd1262: brom_out <= 64'd688271518969994901;
    12'd1263: brom_out <= 64'd6293099328911513541;
    12'd1264: brom_out <= 64'd8022708066944787193;
    12'd1265: brom_out <= 64'd5756412069551489870;
    12'd1266: brom_out <= 64'd3676362487736855076;
    12'd1267: brom_out <= 64'd8145733225084264849;
    12'd1268: brom_out <= 64'd6290626132265462869;
    12'd1269: brom_out <= 64'd3680937565679486776;
    12'd1270: brom_out <= 64'd6506087753855957558;
    12'd1271: brom_out <= 64'd7030390575960316317;
    12'd1272: brom_out <= 64'd710231919379692236;
    12'd1273: brom_out <= 64'd196737007466299716;
    12'd1274: brom_out <= 64'd1613993507937783279;
    12'd1275: brom_out <= 64'd5396535619710247276;
    12'd1276: brom_out <= 64'd3208834222241491524;
    12'd1277: brom_out <= 64'd5426966171602208991;
    12'd1278: brom_out <= 64'd8333424693978152862;
    12'd1279: brom_out <= 64'd8389518664907588327;
    12'd1280: brom_out <= 64'd3843729905249091225;
    12'd1281: brom_out <= 64'd7556005083705865018;
    12'd1282: brom_out <= 64'd4878912351183739034;
    12'd1283: brom_out <= 64'd1333223997973402547;
    12'd1284: brom_out <= 64'd4499316437729491950;
    12'd1285: brom_out <= 64'd166284095181747720;
    12'd1286: brom_out <= 64'd6366904626277906997;
    12'd1287: brom_out <= 64'd586940494231743755;
    12'd1288: brom_out <= 64'd2124775930866948658;
    12'd1289: brom_out <= 64'd1934097126200992158;
    12'd1290: brom_out <= 64'd4446777445590067722;
    12'd1291: brom_out <= 64'd1009392566066621240;
    12'd1292: brom_out <= 64'd5031955862462893125;
    12'd1293: brom_out <= 64'd7906792694894978237;
    12'd1294: brom_out <= 64'd7346123643397775154;
    12'd1295: brom_out <= 64'd8287665031610589475;
    12'd1296: brom_out <= 64'd8597644118437593047;
    12'd1297: brom_out <= 64'd392229208402201833;
    12'd1298: brom_out <= 64'd2996198017684397473;
    12'd1299: brom_out <= 64'd7849377421420064578;
    12'd1300: brom_out <= 64'd1322077954161935913;
    12'd1301: brom_out <= 64'd1736720476753951439;
    12'd1302: brom_out <= 64'd7461692640222935420;
    12'd1303: brom_out <= 64'd330771392035517163;
    12'd1304: brom_out <= 64'd6354329292015303361;
    12'd1305: brom_out <= 64'd3890164895378234331;
    12'd1306: brom_out <= 64'd8222878809597452782;
    12'd1307: brom_out <= 64'd2210258167203109148;
    12'd1308: brom_out <= 64'd5616442847621039958;
    12'd1309: brom_out <= 64'd1981907441775399123;
    12'd1310: brom_out <= 64'd4425836144919842661;
    12'd1311: brom_out <= 64'd3088046495030321430;
    12'd1312: brom_out <= 64'd1103810256172461273;
    12'd1313: brom_out <= 64'd9198512508640536753;
    12'd1314: brom_out <= 64'd8863652633840617892;
    12'd1315: brom_out <= 64'd3811497093829914947;
    12'd1316: brom_out <= 64'd5185697590161398078;
    12'd1317: brom_out <= 64'd2478477691263246336;
    12'd1318: brom_out <= 64'd9041703530576244245;
    12'd1319: brom_out <= 64'd7630500404892957606;
    12'd1320: brom_out <= 64'd2808768542836739127;
    12'd1321: brom_out <= 64'd8506876570223798909;
    12'd1322: brom_out <= 64'd3515447309748454700;
    12'd1323: brom_out <= 64'd5584181301675612560;
    12'd1324: brom_out <= 64'd8076854248606482640;
    12'd1325: brom_out <= 64'd464762712416825453;
    12'd1326: brom_out <= 64'd1212934680674932171;
    12'd1327: brom_out <= 64'd6822705681720740975;
    12'd1328: brom_out <= 64'd1616415171056121951;
    12'd1329: brom_out <= 64'd1858244221136017157;
    12'd1330: brom_out <= 64'd5827250561241730507;
    12'd1331: brom_out <= 64'd344400738107596023;
    12'd1332: brom_out <= 64'd1764465672678590335;
    12'd1333: brom_out <= 64'd5703781165619639802;
    12'd1334: brom_out <= 64'd7628029483406556039;
    12'd1335: brom_out <= 64'd3427262358653674690;
    12'd1336: brom_out <= 64'd2554628785776186101;
    12'd1337: brom_out <= 64'd7220928449331731964;
    12'd1338: brom_out <= 64'd6073433051176488437;
    12'd1339: brom_out <= 64'd1675796553890763688;
    12'd1340: brom_out <= 64'd6274269344659241202;
    12'd1341: brom_out <= 64'd3239268158919342920;
    12'd1342: brom_out <= 64'd857257993458705591;
    12'd1343: brom_out <= 64'd8027273317913045334;
    12'd1344: brom_out <= 64'd7760096502744668708;
    12'd1345: brom_out <= 64'd6293371826854438675;
    12'd1346: brom_out <= 64'd2664415077131265526;
    12'd1347: brom_out <= 64'd6008070311175945680;
    12'd1348: brom_out <= 64'd7774041485289560934;
    12'd1349: brom_out <= 64'd2158497848787983836;
    12'd1350: brom_out <= 64'd7804415236345099072;
    12'd1351: brom_out <= 64'd7766697199279911580;
    12'd1352: brom_out <= 64'd3444196253661916107;
    12'd1353: brom_out <= 64'd7333098404852221282;
    12'd1354: brom_out <= 64'd1408354985644544297;
    12'd1355: brom_out <= 64'd3696418947871042363;
    12'd1356: brom_out <= 64'd4199856302268999704;
    12'd1357: brom_out <= 64'd8667550626171542063;
    12'd1358: brom_out <= 64'd4821450906140543866;
    12'd1359: brom_out <= 64'd5280375575531834917;
    12'd1360: brom_out <= 64'd4742976528600107296;
    12'd1361: brom_out <= 64'd7971062668178884619;
    12'd1362: brom_out <= 64'd2624241653356493808;
    12'd1363: brom_out <= 64'd2943196258777315248;
    12'd1364: brom_out <= 64'd1459241221732760376;
    12'd1365: brom_out <= 64'd3141892699607285042;
    12'd1366: brom_out <= 64'd6779863717923106188;
    12'd1367: brom_out <= 64'd2290981532627662977;
    12'd1368: brom_out <= 64'd2596338163869140878;
    12'd1369: brom_out <= 64'd6132164137524698293;
    12'd1370: brom_out <= 64'd2806704808466864642;
    12'd1371: brom_out <= 64'd1231316600362524550;
    12'd1372: brom_out <= 64'd4878604162374060394;
    12'd1373: brom_out <= 64'd6153996695725736706;
    12'd1374: brom_out <= 64'd8392369886176695753;
    12'd1375: brom_out <= 64'd7381481651865989698;
    12'd1376: brom_out <= 64'd3956250839820662012;
    12'd1377: brom_out <= 64'd4440155139934687816;
    12'd1378: brom_out <= 64'd3410526233184475385;
    12'd1379: brom_out <= 64'd2915613055628798760;
    12'd1380: brom_out <= 64'd3741551785277411008;
    12'd1381: brom_out <= 64'd4095066806824966641;
    12'd1382: brom_out <= 64'd6396076356706250734;
    12'd1383: brom_out <= 64'd6144284829132834422;
    12'd1384: brom_out <= 64'd359462425852779964;
    12'd1385: brom_out <= 64'd2581914814665931179;
    12'd1386: brom_out <= 64'd5164305657351049013;
    12'd1387: brom_out <= 64'd6642437784128992902;
    12'd1388: brom_out <= 64'd7109225250325427391;
    12'd1389: brom_out <= 64'd5881288971893723570;
    12'd1390: brom_out <= 64'd5439199440553482972;
    12'd1391: brom_out <= 64'd8411606107586220522;
    12'd1392: brom_out <= 64'd8842309920213777422;
    12'd1393: brom_out <= 64'd2054983379813627592;
    12'd1394: brom_out <= 64'd3290781571874907490;
    12'd1395: brom_out <= 64'd3450300767690318983;
    12'd1396: brom_out <= 64'd3498405541614573677;
    12'd1397: brom_out <= 64'd7443993893567332439;
    12'd1398: brom_out <= 64'd6785899613309730809;
    12'd1399: brom_out <= 64'd959708987379827311;
    12'd1400: brom_out <= 64'd7756449588084361090;
    12'd1401: brom_out <= 64'd4378670015744532545;
    12'd1402: brom_out <= 64'd7638018630422522758;
    12'd1403: brom_out <= 64'd5513943317299056632;
    12'd1404: brom_out <= 64'd7021500185955960993;
    12'd1405: brom_out <= 64'd3883430424181642244;
    12'd1406: brom_out <= 64'd6441046237530661408;
    12'd1407: brom_out <= 64'd4615964652737150867;
    12'd1408: brom_out <= 64'd953672148357239882;
    12'd1409: brom_out <= 64'd850129065329897070;
    12'd1410: brom_out <= 64'd6867536447291324630;
    12'd1411: brom_out <= 64'd5338739010407762928;
    12'd1412: brom_out <= 64'd4487508645819054224;
    12'd1413: brom_out <= 64'd6655809630869496375;
    12'd1414: brom_out <= 64'd3560640136243016745;
    12'd1415: brom_out <= 64'd2586800327873423869;
    12'd1416: brom_out <= 64'd7881133695797688301;
    12'd1417: brom_out <= 64'd6939558012044222620;
    12'd1418: brom_out <= 64'd8296166227971292689;
    12'd1419: brom_out <= 64'd2809488325196303122;
    12'd1420: brom_out <= 64'd8094583652892052949;
    12'd1421: brom_out <= 64'd3765812450421358809;
    12'd1422: brom_out <= 64'd6661553702290924851;
    12'd1423: brom_out <= 64'd8456238973083966825;
    12'd1424: brom_out <= 64'd2021487688528006903;
    12'd1425: brom_out <= 64'd176821124719014857;
    12'd1426: brom_out <= 64'd2601479532876804086;
    12'd1427: brom_out <= 64'd3102810669834941357;
    12'd1428: brom_out <= 64'd2856594089171996563;
    12'd1429: brom_out <= 64'd1760667119417696491;
    12'd1430: brom_out <= 64'd4727177425397781733;
    12'd1431: brom_out <= 64'd3380819559153913571;
    12'd1432: brom_out <= 64'd7895456088394432312;
    12'd1433: brom_out <= 64'd1813734445697875842;
    12'd1434: brom_out <= 64'd6206618949097304040;
    12'd1435: brom_out <= 64'd5650920825046544428;
    12'd1436: brom_out <= 64'd7655220296250182295;
    12'd1437: brom_out <= 64'd7544241347745579320;
    12'd1438: brom_out <= 64'd727549704694688894;
    12'd1439: brom_out <= 64'd1566328877329519572;
    12'd1440: brom_out <= 64'd3600223915184093972;
    12'd1441: brom_out <= 64'd6135318313250553096;
    12'd1442: brom_out <= 64'd132349231880792967;
    12'd1443: brom_out <= 64'd231521853003109347;
    12'd1444: brom_out <= 64'd8079743228639382862;
    12'd1445: brom_out <= 64'd6017979743130723506;
    12'd1446: brom_out <= 64'd7906606231102725904;
    12'd1447: brom_out <= 64'd703240658030183136;
    12'd1448: brom_out <= 64'd8202248938719511892;
    12'd1449: brom_out <= 64'd5621135452732475537;
    12'd1450: brom_out <= 64'd1440436752413340717;
    12'd1451: brom_out <= 64'd9186394120520577013;
    12'd1452: brom_out <= 64'd1815902719205333795;
    12'd1453: brom_out <= 64'd1156890325131340717;
    12'd1454: brom_out <= 64'd510250283286762805;
    12'd1455: brom_out <= 64'd7003793697811322955;
    12'd1456: brom_out <= 64'd1367942777365248130;
    12'd1457: brom_out <= 64'd8435760018173686736;
    12'd1458: brom_out <= 64'd2294766590646468670;
    12'd1459: brom_out <= 64'd3095476658074671006;
    12'd1460: brom_out <= 64'd459816473559117541;
    12'd1461: brom_out <= 64'd796266968581397676;
    12'd1462: brom_out <= 64'd1609218039696710184;
    12'd1463: brom_out <= 64'd2759828944335218891;
    12'd1464: brom_out <= 64'd3468868502229043904;
    12'd1465: brom_out <= 64'd9046305768736116649;
    12'd1466: brom_out <= 64'd7978421110098049193;
    12'd1467: brom_out <= 64'd902543247035843629;
    12'd1468: brom_out <= 64'd6209991961353846078;
    12'd1469: brom_out <= 64'd7043943473936993612;
    12'd1470: brom_out <= 64'd3718407247601793104;
    12'd1471: brom_out <= 64'd3931580345959350472;
    12'd1472: brom_out <= 64'd6083901335903595160;
    12'd1473: brom_out <= 64'd6824664332907535647;
    12'd1474: brom_out <= 64'd1684476880976375799;
    12'd1475: brom_out <= 64'd8353748286838335736;
    12'd1476: brom_out <= 64'd3101660921827448763;
    12'd1477: brom_out <= 64'd4676099432048506185;
    12'd1478: brom_out <= 64'd353854522259754772;
    12'd1479: brom_out <= 64'd5411283359490134200;
    12'd1480: brom_out <= 64'd3415698136892615027;
    12'd1481: brom_out <= 64'd7966854439247032166;
    12'd1482: brom_out <= 64'd4173694954568519866;
    12'd1483: brom_out <= 64'd5586515692744092763;
    12'd1484: brom_out <= 64'd3411832143259739766;
    12'd1485: brom_out <= 64'd2321500311361878195;
    12'd1486: brom_out <= 64'd4766150303353805783;
    12'd1487: brom_out <= 64'd4189727577864317025;
    12'd1488: brom_out <= 64'd2120186974104516783;
    12'd1489: brom_out <= 64'd2346054488387599429;
    12'd1490: brom_out <= 64'd5821796730151837077;
    12'd1491: brom_out <= 64'd1369377918869971192;
    12'd1492: brom_out <= 64'd6371903036053498044;
    12'd1493: brom_out <= 64'd7515269066369962567;
    12'd1494: brom_out <= 64'd5335315258324712446;
    12'd1495: brom_out <= 64'd2204454453407876475;
    12'd1496: brom_out <= 64'd3987379548559387482;
    12'd1497: brom_out <= 64'd6905936533129222384;
    12'd1498: brom_out <= 64'd6721409961890157156;
    12'd1499: brom_out <= 64'd2790455898821474261;
    12'd1500: brom_out <= 64'd2745037392700744382;
    12'd1501: brom_out <= 64'd3225199442296255605;
    12'd1502: brom_out <= 64'd8886970487032570325;
    12'd1503: brom_out <= 64'd6684109409847610132;
    12'd1504: brom_out <= 64'd2060688072657154489;
    12'd1505: brom_out <= 64'd7631974959581079008;
    12'd1506: brom_out <= 64'd2444995044459230623;
    12'd1507: brom_out <= 64'd5193199074429100689;
    12'd1508: brom_out <= 64'd2852460360135711509;
    12'd1509: brom_out <= 64'd4035422112286893400;
    12'd1510: brom_out <= 64'd789608684700451415;
    12'd1511: brom_out <= 64'd4057000862583680209;
    12'd1512: brom_out <= 64'd6583150359500196198;
    12'd1513: brom_out <= 64'd7750594867189308663;
    12'd1514: brom_out <= 64'd8709515139927426362;
    12'd1515: brom_out <= 64'd9181066187926391646;
    12'd1516: brom_out <= 64'd1351484717233732473;
    12'd1517: brom_out <= 64'd3411154478318304122;
    12'd1518: brom_out <= 64'd423894166336500447;
    12'd1519: brom_out <= 64'd487501164676342059;
    12'd1520: brom_out <= 64'd3160045223296692649;
    12'd1521: brom_out <= 64'd6876782766010347338;
    12'd1522: brom_out <= 64'd6075328695816030615;
    12'd1523: brom_out <= 64'd5607315581519378807;
    12'd1524: brom_out <= 64'd2171281169681126126;
    12'd1525: brom_out <= 64'd7957132803627280334;
    12'd1526: brom_out <= 64'd5415240570595024209;
    12'd1527: brom_out <= 64'd2795954943581859913;
    12'd1528: brom_out <= 64'd1484286524317179508;
    12'd1529: brom_out <= 64'd3630073746381331890;
    12'd1530: brom_out <= 64'd7868389234956506444;
    12'd1531: brom_out <= 64'd6097958069547450574;
    12'd1532: brom_out <= 64'd2217611238809723830;
    12'd1533: brom_out <= 64'd4978123695878332940;
    12'd1534: brom_out <= 64'd928971682581006270;
    12'd1535: brom_out <= 64'd5061989905722694737;
    12'd1536: brom_out <= 64'd5617791344231802350;
    12'd1537: brom_out <= 64'd3311625959390192246;
    12'd1538: brom_out <= 64'd2799145201384261539;
    12'd1539: brom_out <= 64'd6121717495678153306;
    12'd1540: brom_out <= 64'd9130971152851864320;
    12'd1541: brom_out <= 64'd2169428785439006306;
    12'd1542: brom_out <= 64'd363817006911070633;
    12'd1543: brom_out <= 64'd8077220149289012515;
    12'd1544: brom_out <= 64'd2764199408295378392;
    12'd1545: brom_out <= 64'd4572200790955778880;
    12'd1546: brom_out <= 64'd5153420462376781119;
    12'd1547: brom_out <= 64'd8820164290429074374;
    12'd1548: brom_out <= 64'd6828356927799211956;
    12'd1549: brom_out <= 64'd4928657927327845097;
    12'd1550: brom_out <= 64'd2626402754532212200;
    12'd1551: brom_out <= 64'd957663858492823873;
    12'd1552: brom_out <= 64'd4659108819977211531;
    12'd1553: brom_out <= 64'd4008307678287682078;
    12'd1554: brom_out <= 64'd3630244555345427809;
    12'd1555: brom_out <= 64'd5162240120750053334;
    12'd1556: brom_out <= 64'd5992236777911864655;
    12'd1557: brom_out <= 64'd21240054144111511;
    12'd1558: brom_out <= 64'd8213520103588895170;
    12'd1559: brom_out <= 64'd5886493698929414728;
    12'd1560: brom_out <= 64'd6341707651478976599;
    12'd1561: brom_out <= 64'd7667751154799082802;
    12'd1562: brom_out <= 64'd237652332054158574;
    12'd1563: brom_out <= 64'd8445874054791808278;
    12'd1564: brom_out <= 64'd1116527593943410644;
    12'd1565: brom_out <= 64'd5834422649485691430;
    12'd1566: brom_out <= 64'd2610995018984948356;
    12'd1567: brom_out <= 64'd8992065833585364210;
    12'd1568: brom_out <= 64'd3783999585861312710;
    12'd1569: brom_out <= 64'd8659767712472380210;
    12'd1570: brom_out <= 64'd1451024343543556476;
    12'd1571: brom_out <= 64'd852251189757033736;
    12'd1572: brom_out <= 64'd715272894832880454;
    12'd1573: brom_out <= 64'd3170151885362480463;
    12'd1574: brom_out <= 64'd7963579077243854117;
    12'd1575: brom_out <= 64'd4409479336568326293;
    12'd1576: brom_out <= 64'd8238224820786296794;
    12'd1577: brom_out <= 64'd4476045774402502806;
    12'd1578: brom_out <= 64'd2173707138548862621;
    12'd1579: brom_out <= 64'd6474722828429963680;
    12'd1580: brom_out <= 64'd3534484640152137503;
    12'd1581: brom_out <= 64'd8299199171065342576;
    12'd1582: brom_out <= 64'd4645071257540983012;
    12'd1583: brom_out <= 64'd2271101635375968800;
    12'd1584: brom_out <= 64'd5044931045435287860;
    12'd1585: brom_out <= 64'd1371172093890878646;
    12'd1586: brom_out <= 64'd3421777070366820959;
    12'd1587: brom_out <= 64'd4775821216533904327;
    12'd1588: brom_out <= 64'd6731965169435440516;
    12'd1589: brom_out <= 64'd6240908704213519302;
    12'd1590: brom_out <= 64'd9180299276538237891;
    12'd1591: brom_out <= 64'd3826833899262929350;
    12'd1592: brom_out <= 64'd1358546831763501466;
    12'd1593: brom_out <= 64'd5795760311661694782;
    12'd1594: brom_out <= 64'd857649613222965065;
    12'd1595: brom_out <= 64'd5374038621152501313;
    12'd1596: brom_out <= 64'd1195287042107083358;
    12'd1597: brom_out <= 64'd5814958504459929101;
    12'd1598: brom_out <= 64'd5213930122402843181;
    12'd1599: brom_out <= 64'd3814003116314377089;
    12'd1600: brom_out <= 64'd4360836354755007548;
    12'd1601: brom_out <= 64'd2807089391805868739;
    12'd1602: brom_out <= 64'd5401705995168057573;
    12'd1603: brom_out <= 64'd7565883564426729174;
    12'd1604: brom_out <= 64'd5695113735564493386;
    12'd1605: brom_out <= 64'd973486816132687795;
    12'd1606: brom_out <= 64'd5295305162382387292;
    12'd1607: brom_out <= 64'd7246454730830313036;
    12'd1608: brom_out <= 64'd3338745277371104260;
    12'd1609: brom_out <= 64'd164458380228977682;
    12'd1610: brom_out <= 64'd6611118261441405900;
    12'd1611: brom_out <= 64'd194947333109386454;
    12'd1612: brom_out <= 64'd2856515524884644876;
    12'd1613: brom_out <= 64'd5993844322502066692;
    12'd1614: brom_out <= 64'd4610665961523289949;
    12'd1615: brom_out <= 64'd3613202757720993929;
    12'd1616: brom_out <= 64'd3492678159767424326;
    12'd1617: brom_out <= 64'd1035633680400379250;
    12'd1618: brom_out <= 64'd1107635849814668979;
    12'd1619: brom_out <= 64'd6121644004340863046;
    12'd1620: brom_out <= 64'd4142681969498947811;
    12'd1621: brom_out <= 64'd5106407504416289347;
    12'd1622: brom_out <= 64'd4587503492636103025;
    12'd1623: brom_out <= 64'd1549219934878699976;
    12'd1624: brom_out <= 64'd6112709126884308384;
    12'd1625: brom_out <= 64'd1536559248545772238;
    12'd1626: brom_out <= 64'd4564261353425194389;
    12'd1627: brom_out <= 64'd4407786248107552167;
    12'd1628: brom_out <= 64'd8462729403610917864;
    12'd1629: brom_out <= 64'd7635802621249192949;
    12'd1630: brom_out <= 64'd5617373606608073906;
    12'd1631: brom_out <= 64'd6278949468837188216;
    12'd1632: brom_out <= 64'd4618095554046765688;
    12'd1633: brom_out <= 64'd2001877912459119594;
    12'd1634: brom_out <= 64'd5627259502194020199;
    12'd1635: brom_out <= 64'd6838396562566836729;
    12'd1636: brom_out <= 64'd3093321946376148894;
    12'd1637: brom_out <= 64'd3377148768122421051;
    12'd1638: brom_out <= 64'd2625927586413902378;
    12'd1639: brom_out <= 64'd8720594263944441184;
    12'd1640: brom_out <= 64'd1186120250261651295;
    12'd1641: brom_out <= 64'd8427722037080059434;
    12'd1642: brom_out <= 64'd6160205427239796113;
    12'd1643: brom_out <= 64'd9142186737552927218;
    12'd1644: brom_out <= 64'd8275074185071956353;
    12'd1645: brom_out <= 64'd3643958317708593014;
    12'd1646: brom_out <= 64'd2698627880457448294;
    12'd1647: brom_out <= 64'd3060636953399987899;
    12'd1648: brom_out <= 64'd1670522412820839339;
    12'd1649: brom_out <= 64'd433728210396661704;
    12'd1650: brom_out <= 64'd3192416431815291977;
    12'd1651: brom_out <= 64'd217683746062300453;
    12'd1652: brom_out <= 64'd190138040081956250;
    12'd1653: brom_out <= 64'd6096016772228045947;
    12'd1654: brom_out <= 64'd4890768885230644118;
    12'd1655: brom_out <= 64'd4594351722144035398;
    12'd1656: brom_out <= 64'd1654928964314873373;
    12'd1657: brom_out <= 64'd895906353740599246;
    12'd1658: brom_out <= 64'd697152114074171637;
    12'd1659: brom_out <= 64'd6653468028538889837;
    12'd1660: brom_out <= 64'd7606147805583021835;
    12'd1661: brom_out <= 64'd3154851592447277802;
    12'd1662: brom_out <= 64'd8750950506552978663;
    12'd1663: brom_out <= 64'd6428260343660144231;
    12'd1664: brom_out <= 64'd7110756539493835260;
    12'd1665: brom_out <= 64'd2192138033866419697;
    12'd1666: brom_out <= 64'd7305100591989071130;
    12'd1667: brom_out <= 64'd5735924744281119282;
    12'd1668: brom_out <= 64'd2778425647746173460;
    12'd1669: brom_out <= 64'd5399144814289903092;
    12'd1670: brom_out <= 64'd5344955090064714738;
    12'd1671: brom_out <= 64'd1844186876280008733;
    12'd1672: brom_out <= 64'd3718083491073040252;
    12'd1673: brom_out <= 64'd7698480780335511647;
    12'd1674: brom_out <= 64'd8265472217763378566;
    12'd1675: brom_out <= 64'd7531439844359758975;
    12'd1676: brom_out <= 64'd8171984989099906491;
    12'd1677: brom_out <= 64'd8856053219407297478;
    12'd1678: brom_out <= 64'd8775554507670322674;
    12'd1679: brom_out <= 64'd6541234765908904047;
    12'd1680: brom_out <= 64'd4557700549816687005;
    12'd1681: brom_out <= 64'd2262383647763924369;
    12'd1682: brom_out <= 64'd1242142187437704347;
    12'd1683: brom_out <= 64'd5265272503518076052;
    12'd1684: brom_out <= 64'd3136793583253461037;
    12'd1685: brom_out <= 64'd796967671211981828;
    12'd1686: brom_out <= 64'd7642072530786664933;
    12'd1687: brom_out <= 64'd734856006618963226;
    12'd1688: brom_out <= 64'd221067181956826324;
    12'd1689: brom_out <= 64'd3722433187835893578;
    12'd1690: brom_out <= 64'd6491983198110424931;
    12'd1691: brom_out <= 64'd9082617714353364049;
    12'd1692: brom_out <= 64'd6602110944466075840;
    12'd1693: brom_out <= 64'd1085578947392235392;
    12'd1694: brom_out <= 64'd3616132668740753638;
    12'd1695: brom_out <= 64'd3703896699573254429;
    12'd1696: brom_out <= 64'd2118076072849861137;
    12'd1697: brom_out <= 64'd3043476125592443538;
    12'd1698: brom_out <= 64'd3210435579848204682;
    12'd1699: brom_out <= 64'd8697093929647739149;
    12'd1700: brom_out <= 64'd8841447671122217172;
    12'd1701: brom_out <= 64'd491533638022032998;
    12'd1702: brom_out <= 64'd3144422523795751301;
    12'd1703: brom_out <= 64'd2510322458979468606;
    12'd1704: brom_out <= 64'd108103996902987755;
    12'd1705: brom_out <= 64'd8575727335521542901;
    12'd1706: brom_out <= 64'd5717679017859454353;
    12'd1707: brom_out <= 64'd4041080959967286788;
    12'd1708: brom_out <= 64'd5726899559991123300;
    12'd1709: brom_out <= 64'd789285590662622296;
    12'd1710: brom_out <= 64'd8634143088716469639;
    12'd1711: brom_out <= 64'd4230337959405382367;
    12'd1712: brom_out <= 64'd2959784714975049404;
    12'd1713: brom_out <= 64'd2804864706059028877;
    12'd1714: brom_out <= 64'd4711440369215415820;
    12'd1715: brom_out <= 64'd8861845489832604060;
    12'd1716: brom_out <= 64'd540676285453317412;
    12'd1717: brom_out <= 64'd1236972992005525903;
    12'd1718: brom_out <= 64'd1625756756431133274;
    12'd1719: brom_out <= 64'd8811191242823468048;
    12'd1720: brom_out <= 64'd2182142605934843773;
    12'd1721: brom_out <= 64'd8722561625366557139;
    12'd1722: brom_out <= 64'd2548943407954106725;
    12'd1723: brom_out <= 64'd5445744561058896781;
    12'd1724: brom_out <= 64'd717772132402160768;
    12'd1725: brom_out <= 64'd3890495947032713939;
    12'd1726: brom_out <= 64'd763114800931767035;
    12'd1727: brom_out <= 64'd9139193084538540417;
    12'd1728: brom_out <= 64'd9214823842518320290;
    12'd1729: brom_out <= 64'd7106124249430698532;
    12'd1730: brom_out <= 64'd4356193493955929660;
    12'd1731: brom_out <= 64'd4967125163733076709;
    12'd1732: brom_out <= 64'd10155564005954711;
    12'd1733: brom_out <= 64'd1780292907307957066;
    12'd1734: brom_out <= 64'd3820834095675889318;
    12'd1735: brom_out <= 64'd900808569202260949;
    12'd1736: brom_out <= 64'd6488067714213829364;
    12'd1737: brom_out <= 64'd550889388219269783;
    12'd1738: brom_out <= 64'd8849440942935126123;
    12'd1739: brom_out <= 64'd2186610694973659466;
    12'd1740: brom_out <= 64'd1225871290653235241;
    12'd1741: brom_out <= 64'd361423748258118745;
    12'd1742: brom_out <= 64'd4506876142162943112;
    12'd1743: brom_out <= 64'd2010875364009173480;
    12'd1744: brom_out <= 64'd5129958208395442412;
    12'd1745: brom_out <= 64'd3083099219996215074;
    12'd1746: brom_out <= 64'd8837937225769182693;
    12'd1747: brom_out <= 64'd1146124925862289999;
    12'd1748: brom_out <= 64'd2034031322230827706;
    12'd1749: brom_out <= 64'd1105586051061267328;
    12'd1750: brom_out <= 64'd3714772894063112217;
    12'd1751: brom_out <= 64'd2167058803693745213;
    12'd1752: brom_out <= 64'd2721304064985168695;
    12'd1753: brom_out <= 64'd8591940083993862567;
    12'd1754: brom_out <= 64'd2460648692420495320;
    12'd1755: brom_out <= 64'd2508975431031940143;
    12'd1756: brom_out <= 64'd2268060123631796342;
    12'd1757: brom_out <= 64'd5900959382402831706;
    12'd1758: brom_out <= 64'd4277461058176170045;
    12'd1759: brom_out <= 64'd7184971508331829241;
    12'd1760: brom_out <= 64'd43318055585353588;
    12'd1761: brom_out <= 64'd6296341197324853931;
    12'd1762: brom_out <= 64'd3632225739685008221;
    12'd1763: brom_out <= 64'd1937376737223836732;
    12'd1764: brom_out <= 64'd8891709454381057004;
    12'd1765: brom_out <= 64'd6012706981821976828;
    12'd1766: brom_out <= 64'd8109043667728856577;
    12'd1767: brom_out <= 64'd3278792716225804354;
    12'd1768: brom_out <= 64'd2423438989550509849;
    12'd1769: brom_out <= 64'd7191337575891006538;
    12'd1770: brom_out <= 64'd3385836186374320930;
    12'd1771: brom_out <= 64'd3269245869410515417;
    12'd1772: brom_out <= 64'd7117238200784564383;
    12'd1773: brom_out <= 64'd5499757955899089860;
    12'd1774: brom_out <= 64'd959531988668586204;
    12'd1775: brom_out <= 64'd4776210228079752720;
    12'd1776: brom_out <= 64'd9118542527250028416;
    12'd1777: brom_out <= 64'd4267248588058011112;
    12'd1778: brom_out <= 64'd3249971412615813818;
    12'd1779: brom_out <= 64'd161549653327374463;
    12'd1780: brom_out <= 64'd8052839275297477171;
    12'd1781: brom_out <= 64'd2715847114076104891;
    12'd1782: brom_out <= 64'd9135596727390081326;
    12'd1783: brom_out <= 64'd3216942250772631953;
    12'd1784: brom_out <= 64'd942648120926805071;
    12'd1785: brom_out <= 64'd8873623029041645127;
    12'd1786: brom_out <= 64'd6839157252365283657;
    12'd1787: brom_out <= 64'd8320995123289679476;
    12'd1788: brom_out <= 64'd3118176081677087950;
    12'd1789: brom_out <= 64'd351009294231000662;
    12'd1790: brom_out <= 64'd7272488507232229518;
    12'd1791: brom_out <= 64'd7629084228617682799;
    12'd1792: brom_out <= 64'd7799879935344187323;
    12'd1793: brom_out <= 64'd2449120746788553391;
    12'd1794: brom_out <= 64'd2272934008799617957;
    12'd1795: brom_out <= 64'd7303112304720635750;
    12'd1796: brom_out <= 64'd760300682967404465;
    12'd1797: brom_out <= 64'd1402256476136217707;
    12'd1798: brom_out <= 64'd3391459215294077910;
    12'd1799: brom_out <= 64'd4259947076671469396;
    12'd1800: brom_out <= 64'd5451374971511350464;
    12'd1801: brom_out <= 64'd8462210498215899141;
    12'd1802: brom_out <= 64'd9082017356295096735;
    12'd1803: brom_out <= 64'd1802003130975063954;
    12'd1804: brom_out <= 64'd8272790162005470148;
    12'd1805: brom_out <= 64'd6423625592867496534;
    12'd1806: brom_out <= 64'd8732913552528363436;
    12'd1807: brom_out <= 64'd7670081967714960325;
    12'd1808: brom_out <= 64'd5788755231736737505;
    12'd1809: brom_out <= 64'd2241205217165107414;
    12'd1810: brom_out <= 64'd7557464083934741533;
    12'd1811: brom_out <= 64'd5680215377256052946;
    12'd1812: brom_out <= 64'd4742551049497877389;
    12'd1813: brom_out <= 64'd3915421441849566989;
    12'd1814: brom_out <= 64'd4419464548329866583;
    12'd1815: brom_out <= 64'd2269193766469671833;
    12'd1816: brom_out <= 64'd125145389407238227;
    12'd1817: brom_out <= 64'd4322543213393404369;
    12'd1818: brom_out <= 64'd1730084178090489027;
    12'd1819: brom_out <= 64'd6418502706900467582;
    12'd1820: brom_out <= 64'd5486407041020905443;
    12'd1821: brom_out <= 64'd6893095921796554469;
    12'd1822: brom_out <= 64'd1276085309250879688;
    12'd1823: brom_out <= 64'd8136986804572815553;
    12'd1824: brom_out <= 64'd8878014989630440906;
    12'd1825: brom_out <= 64'd2054499947427697277;
    12'd1826: brom_out <= 64'd4958364417677015727;
    12'd1827: brom_out <= 64'd8639883397318540390;
    12'd1828: brom_out <= 64'd6405046534155161981;
    12'd1829: brom_out <= 64'd3855991029263222897;
    12'd1830: brom_out <= 64'd3849863099847043327;
    12'd1831: brom_out <= 64'd5461834086845665801;
    12'd1832: brom_out <= 64'd5383822019583725910;
    12'd1833: brom_out <= 64'd6843674835657216928;
    12'd1834: brom_out <= 64'd8817907421746805699;
    12'd1835: brom_out <= 64'd1310096281335176417;
    12'd1836: brom_out <= 64'd1591164740821625308;
    12'd1837: brom_out <= 64'd1130529612131441025;
    12'd1838: brom_out <= 64'd1901563757671036646;
    12'd1839: brom_out <= 64'd5904894196451122007;
    12'd1840: brom_out <= 64'd3516589675860114141;
    12'd1841: brom_out <= 64'd6417488381876655358;
    12'd1842: brom_out <= 64'd8273432024380977131;
    12'd1843: brom_out <= 64'd7290240891834356013;
    12'd1844: brom_out <= 64'd5019962465176564987;
    12'd1845: brom_out <= 64'd3690342459317836959;
    12'd1846: brom_out <= 64'd8304681131298863243;
    12'd1847: brom_out <= 64'd46919950701852262;
    12'd1848: brom_out <= 64'd1600285536644558808;
    12'd1849: brom_out <= 64'd2945395305975380311;
    12'd1850: brom_out <= 64'd5916834261026815385;
    12'd1851: brom_out <= 64'd340320363819378969;
    12'd1852: brom_out <= 64'd7836292489991860779;
    12'd1853: brom_out <= 64'd1653685435908513775;
    12'd1854: brom_out <= 64'd6280676770146501670;
    12'd1855: brom_out <= 64'd8879135449218147244;
    12'd1856: brom_out <= 64'd6482325237945511459;
    12'd1857: brom_out <= 64'd3499913247207209486;
    12'd1858: brom_out <= 64'd267529195173947995;
    12'd1859: brom_out <= 64'd7095245265796401803;
    12'd1860: brom_out <= 64'd6167588276897908036;
    12'd1861: brom_out <= 64'd4995587661985367569;
    12'd1862: brom_out <= 64'd8847788509959360291;
    12'd1863: brom_out <= 64'd5379019455004121810;
    12'd1864: brom_out <= 64'd721609409607618860;
    12'd1865: brom_out <= 64'd346852958683529622;
    12'd1866: brom_out <= 64'd5375083910833564937;
    12'd1867: brom_out <= 64'd5545978348244844247;
    12'd1868: brom_out <= 64'd8328070745302195818;
    12'd1869: brom_out <= 64'd7352408759901583521;
    12'd1870: brom_out <= 64'd4025627965310674316;
    12'd1871: brom_out <= 64'd2601171251875055375;
    12'd1872: brom_out <= 64'd2048422362597070268;
    12'd1873: brom_out <= 64'd8698121772985835948;
    12'd1874: brom_out <= 64'd3935113794159243174;
    12'd1875: brom_out <= 64'd4934207483627279877;
    12'd1876: brom_out <= 64'd3392029771587990390;
    12'd1877: brom_out <= 64'd8272834808806498581;
    12'd1878: brom_out <= 64'd2758558891568233325;
    12'd1879: brom_out <= 64'd6047100775382455619;
    12'd1880: brom_out <= 64'd1144709855391150131;
    12'd1881: brom_out <= 64'd1322622329280553132;
    12'd1882: brom_out <= 64'd6373914377105343036;
    12'd1883: brom_out <= 64'd6780464550986213562;
    12'd1884: brom_out <= 64'd8205443440992883590;
    12'd1885: brom_out <= 64'd5432062150452453140;
    12'd1886: brom_out <= 64'd8563341485109490608;
    12'd1887: brom_out <= 64'd6344884790361459878;
    12'd1888: brom_out <= 64'd6491230813524270104;
    12'd1889: brom_out <= 64'd5146189575352380294;
    12'd1890: brom_out <= 64'd5050731834744131339;
    12'd1891: brom_out <= 64'd6978185229619619995;
    12'd1892: brom_out <= 64'd8914416700219747609;
    12'd1893: brom_out <= 64'd6507729040352245500;
    12'd1894: brom_out <= 64'd7348421852782387132;
    12'd1895: brom_out <= 64'd25048117730675259;
    12'd1896: brom_out <= 64'd5471072111151109148;
    12'd1897: brom_out <= 64'd2592674720440310106;
    12'd1898: brom_out <= 64'd8590512243527039086;
    12'd1899: brom_out <= 64'd128308396099142330;
    12'd1900: brom_out <= 64'd6468727959095527758;
    12'd1901: brom_out <= 64'd8619483919931264003;
    12'd1902: brom_out <= 64'd1795515970786001141;
    12'd1903: brom_out <= 64'd348664825324288597;
    12'd1904: brom_out <= 64'd2974750146664762930;
    12'd1905: brom_out <= 64'd4270523319905305484;
    12'd1906: brom_out <= 64'd6008836189323739193;
    12'd1907: brom_out <= 64'd1166127705953489199;
    12'd1908: brom_out <= 64'd1654167995963963661;
    12'd1909: brom_out <= 64'd8690366304852788805;
    12'd1910: brom_out <= 64'd3619470125316298575;
    12'd1911: brom_out <= 64'd1841710140923991090;
    12'd1912: brom_out <= 64'd2890183973319040277;
    12'd1913: brom_out <= 64'd2331110739161486355;
    12'd1914: brom_out <= 64'd5119555131095889488;
    12'd1915: brom_out <= 64'd3449673358908680369;
    12'd1916: brom_out <= 64'd8963269062908814356;
    12'd1917: brom_out <= 64'd4361885023796029498;
    12'd1918: brom_out <= 64'd7616945085266707101;
    12'd1919: brom_out <= 64'd106484800563207163;
    12'd1920: brom_out <= 64'd152972107828962887;
    12'd1921: brom_out <= 64'd2771557478354280102;
    12'd1922: brom_out <= 64'd626085302192577848;
    12'd1923: brom_out <= 64'd4979779557253162501;
    12'd1924: brom_out <= 64'd1292738030668931808;
    12'd1925: brom_out <= 64'd330367904191560310;
    12'd1926: brom_out <= 64'd2127672530715019873;
    12'd1927: brom_out <= 64'd5949769470116563528;
    12'd1928: brom_out <= 64'd1162314052316656334;
    12'd1929: brom_out <= 64'd8497157738710866554;
    12'd1930: brom_out <= 64'd5784014104914335116;
    12'd1931: brom_out <= 64'd1431546682450061430;
    12'd1932: brom_out <= 64'd620672310144596356;
    12'd1933: brom_out <= 64'd6906723235701454772;
    12'd1934: brom_out <= 64'd441445969502826770;
    12'd1935: brom_out <= 64'd7280976441114932219;
    12'd1936: brom_out <= 64'd7656385359106811055;
    12'd1937: brom_out <= 64'd1941454423349872774;
    12'd1938: brom_out <= 64'd3350475165838631035;
    12'd1939: brom_out <= 64'd8883676960518262680;
    12'd1940: brom_out <= 64'd6098642081478079379;
    12'd1941: brom_out <= 64'd6880083817266214666;
    12'd1942: brom_out <= 64'd1833072023934069218;
    12'd1943: brom_out <= 64'd7491702495939745603;
    12'd1944: brom_out <= 64'd4317082530005278608;
    12'd1945: brom_out <= 64'd8937159405096425696;
    12'd1946: brom_out <= 64'd921007660662007758;
    12'd1947: brom_out <= 64'd2266398681594291791;
    12'd1948: brom_out <= 64'd2054367836150137383;
    12'd1949: brom_out <= 64'd7038018752512707129;
    12'd1950: brom_out <= 64'd3752104441186131359;
    12'd1951: brom_out <= 64'd2132856335439328310;
    12'd1952: brom_out <= 64'd7169216581217846864;
    12'd1953: brom_out <= 64'd3268163730688804694;
    12'd1954: brom_out <= 64'd1367202631222351884;
    12'd1955: brom_out <= 64'd6326853994154594052;
    12'd1956: brom_out <= 64'd7006492825336182042;
    12'd1957: brom_out <= 64'd3067417224551825324;
    12'd1958: brom_out <= 64'd8390289897894421784;
    12'd1959: brom_out <= 64'd6459981822124125414;
    12'd1960: brom_out <= 64'd3968889466496500974;
    12'd1961: brom_out <= 64'd8313419918288321449;
    12'd1962: brom_out <= 64'd3902232027484765702;
    12'd1963: brom_out <= 64'd7654783203964713034;
    12'd1964: brom_out <= 64'd8643208206667495248;
    12'd1965: brom_out <= 64'd7525524187409032073;
    12'd1966: brom_out <= 64'd2596774662051353996;
    12'd1967: brom_out <= 64'd4684897218052723440;
    12'd1968: brom_out <= 64'd7265808700877099470;
    12'd1969: brom_out <= 64'd5487416088241385428;
    12'd1970: brom_out <= 64'd5547609792552593689;
    12'd1971: brom_out <= 64'd5593793850381701264;
    12'd1972: brom_out <= 64'd2597346571447091066;
    12'd1973: brom_out <= 64'd4521586504942949225;
    12'd1974: brom_out <= 64'd5951244987899276014;
    12'd1975: brom_out <= 64'd545189652856346927;
    12'd1976: brom_out <= 64'd3342289812197437073;
    12'd1977: brom_out <= 64'd3863895514183921091;
    12'd1978: brom_out <= 64'd620228462665540912;
    12'd1979: brom_out <= 64'd7837777609722958241;
    12'd1980: brom_out <= 64'd530449859038129497;
    12'd1981: brom_out <= 64'd5231823286612848958;
    12'd1982: brom_out <= 64'd6989069606975543519;
    12'd1983: brom_out <= 64'd8440189420678092499;
    12'd1984: brom_out <= 64'd8802530656487450100;
    12'd1985: brom_out <= 64'd5957182057853295242;
    12'd1986: brom_out <= 64'd5651925408707418368;
    12'd1987: brom_out <= 64'd7170299547819584987;
    12'd1988: brom_out <= 64'd5760921106279527014;
    12'd1989: brom_out <= 64'd8774930317025118813;
    12'd1990: brom_out <= 64'd2514994721960832184;
    12'd1991: brom_out <= 64'd8156350698089245497;
    12'd1992: brom_out <= 64'd8092028202770013595;
    12'd1993: brom_out <= 64'd2945051867074066815;
    12'd1994: brom_out <= 64'd3048107258014773416;
    12'd1995: brom_out <= 64'd5287276224121412201;
    12'd1996: brom_out <= 64'd1977473528172302974;
    12'd1997: brom_out <= 64'd837914530468971941;
    12'd1998: brom_out <= 64'd86028093078837575;
    12'd1999: brom_out <= 64'd7178987986310357994;
    12'd2000: brom_out <= 64'd2833080917595641053;
    12'd2001: brom_out <= 64'd4850396737100695623;
    12'd2002: brom_out <= 64'd730707792149410394;
    12'd2003: brom_out <= 64'd5837938833226886992;
    12'd2004: brom_out <= 64'd3220167084924640416;
    12'd2005: brom_out <= 64'd1137030056806412582;
    12'd2006: brom_out <= 64'd8764961600979841729;
    12'd2007: brom_out <= 64'd6982180111368799950;
    12'd2008: brom_out <= 64'd4230367111019978792;
    12'd2009: brom_out <= 64'd8472744867647843428;
    12'd2010: brom_out <= 64'd6781316032784920429;
    12'd2011: brom_out <= 64'd7303621341712018276;
    12'd2012: brom_out <= 64'd8700037870304188663;
    12'd2013: brom_out <= 64'd7576665871445803703;
    12'd2014: brom_out <= 64'd3153589616895710680;
    12'd2015: brom_out <= 64'd6926179402678303735;
    12'd2016: brom_out <= 64'd5649029047297330701;
    12'd2017: brom_out <= 64'd2699505448424011853;
    12'd2018: brom_out <= 64'd4753479972855109987;
    12'd2019: brom_out <= 64'd4042493884873251407;
    12'd2020: brom_out <= 64'd7461760175322938184;
    12'd2021: brom_out <= 64'd7925326134315901832;
    12'd2022: brom_out <= 64'd4556779578756386008;
    12'd2023: brom_out <= 64'd1234392369493637338;
    12'd2024: brom_out <= 64'd948434792261929775;
    12'd2025: brom_out <= 64'd3596222308311112711;
    12'd2026: brom_out <= 64'd7267305599223558729;
    12'd2027: brom_out <= 64'd8337173169099121667;
    12'd2028: brom_out <= 64'd7989457675622623999;
    12'd2029: brom_out <= 64'd1673908163281639090;
    12'd2030: brom_out <= 64'd7773356441300667323;
    12'd2031: brom_out <= 64'd729021657513626886;
    12'd2032: brom_out <= 64'd2365490612534447454;
    12'd2033: brom_out <= 64'd511190818015486693;
    12'd2034: brom_out <= 64'd5151352955011766623;
    12'd2035: brom_out <= 64'd6911759165101450306;
    12'd2036: brom_out <= 64'd7034322664781632447;
    12'd2037: brom_out <= 64'd1506390817673699154;
    12'd2038: brom_out <= 64'd4632150496265362581;
    12'd2039: brom_out <= 64'd7056931086227913840;
    12'd2040: brom_out <= 64'd6665507664676739661;
    12'd2041: brom_out <= 64'd2341354910130103652;
    12'd2042: brom_out <= 64'd8477174779707217963;
    12'd2043: brom_out <= 64'd5491683881414165578;
    12'd2044: brom_out <= 64'd1868094419334665511;
    12'd2045: brom_out <= 64'd5881135019807506724;
    12'd2046: brom_out <= 64'd3013299072814627077;
    12'd2047: brom_out <= 64'd6099799931271616695;
    default: brom_out <= 64'h1;
    endcase
end

generate
    if(DELAY == 1) begin
        assign b = brom_out;
    end
endgenerate

endmodule

