`timescale 1ns / 1ps

//-------------------------------------------------------------------------------------------------

module tw_rom_1
#(
    parameter LOGN  = 1,
    parameter LOGQ  = 64,
    parameter DELAY = 1,
    parameter STAGE = 1
)(
    input            clk,
    input [LOGN-1:0] raddr,
    output[LOGQ-1:0] b
);

(* rom_style = "distributed" *)
reg [LOGQ-1:0] brom_out, brom_out2;

always @(posedge clk) begin
    case(raddr[STAGE-1:0])
    2'd0: brom_out <= 64'd9223372036854251519;
    2'd1: brom_out <= 64'd6551015095526749063;
    default: brom_out <= 64'h1;
    endcase
end

generate
    if(DELAY == 1) begin
        assign b = brom_out;
    end
endgenerate

endmodule

//-------------------------------------------------------------------------------------------------

module tw_rom_2
#(
    parameter LOGN  = 2,
    parameter LOGQ  = 64,
    parameter DELAY = 1,
    parameter STAGE = 1
)(
    input            clk,
    input [LOGN-1:0] raddr,
    output[LOGQ-1:0] b
);

(* rom_style = "distributed" *)
reg [LOGQ-1:0] brom_out, brom_out2;

always @(posedge clk) begin
    case(raddr[STAGE-1:0])
    3'd0: brom_out <= 64'd9223372036854251519;
    3'd1: brom_out <= 64'd5976068779477487504;
    3'd2: brom_out <= 64'd6551015095526749063;
    3'd3: brom_out <= 64'd3392617565049336557;
    default: brom_out <= 64'h1;
    endcase
end

generate
    if(DELAY == 1) begin
        assign b = brom_out;
    end
endgenerate

endmodule

//-------------------------------------------------------------------------------------------------

module tw_rom_3
#(
    parameter LOGN  = 3,
    parameter LOGQ  = 64,
    parameter DELAY = 1,
    parameter STAGE = 1
)(
    input            clk,
    input [LOGN-1:0] raddr,
    output[LOGQ-1:0] b
);

(* rom_style = "distributed" *)
reg [LOGQ-1:0] brom_out, brom_out2;

always @(posedge clk) begin
    case(raddr[STAGE-1:0])
    4'd0: brom_out <= 64'd9223372036854251519;
    4'd1: brom_out <= 64'd2881966912403406253;
    4'd2: brom_out <= 64'd5976068779477487504;
    4'd3: brom_out <= 64'd5792979130194094298;
    4'd4: brom_out <= 64'd6551015095526749063;
    4'd5: brom_out <= 64'd2991444385089030097;
    4'd6: brom_out <= 64'd3392617565049336557;
    4'd7: brom_out <= 64'd699101306064864663;
    default: brom_out <= 64'h1;
    endcase
end

generate
    if(DELAY == 1) begin
        assign b = brom_out;
    end
endgenerate

endmodule

//-------------------------------------------------------------------------------------------------

module tw_rom_4
#(
    parameter LOGN  = 4,
    parameter LOGQ  = 64,
    parameter DELAY = 1,
    parameter STAGE = 1
)(
    input            clk,
    input [LOGN-1:0] raddr,
    output[LOGQ-1:0] b
);

(* rom_style = "distributed" *)
reg [LOGQ-1:0] brom_out, brom_out2;

always @(posedge clk) begin
    case(raddr[STAGE-1:0])
    5'd0: brom_out <= 64'd9223372036854251519;
    5'd1: brom_out <= 64'd5917339183240377480;
    5'd2: brom_out <= 64'd2881966912403406253;
    5'd3: brom_out <= 64'd7147821265559899415;
    5'd4: brom_out <= 64'd5976068779477487504;
    5'd5: brom_out <= 64'd4066724171054462909;
    5'd6: brom_out <= 64'd5792979130194094298;
    5'd7: brom_out <= 64'd2803267708398697040;
    5'd8: brom_out <= 64'd6551015095526749063;
    5'd9: brom_out <= 64'd5908178380096272369;
    5'd10: brom_out <= 64'd2991444385089030097;
    5'd11: brom_out <= 64'd7646914504675205489;
    5'd12: brom_out <= 64'd3392617565049336557;
    5'd13: brom_out <= 64'd1002059954001900696;
    5'd14: brom_out <= 64'd699101306064864663;
    5'd15: brom_out <= 64'd1670791095363685175;
    default: brom_out <= 64'h1;
    endcase
end

generate
    if(DELAY == 1) begin
        assign b = brom_out;
    end
endgenerate

endmodule

//-------------------------------------------------------------------------------------------------

module tw_rom_5
#(
    parameter LOGN  = 5,
    parameter LOGQ  = 64,
    parameter DELAY = 1,
    parameter STAGE = 1
)(
    input            clk,
    input [LOGN-1:0] raddr,
    output[LOGQ-1:0] b
);

(* rom_style = "distributed" *)
reg [LOGQ-1:0] brom_out, brom_out2;

always @(posedge clk) begin
    case(raddr[STAGE-1:0])
    6'd0: brom_out <= 64'd9223372036854251519;
    6'd1: brom_out <= 64'd8706294438413809553;
    6'd2: brom_out <= 64'd5917339183240377480;
    6'd3: brom_out <= 64'd4110363107264655732;
    6'd4: brom_out <= 64'd2881966912403406253;
    6'd5: brom_out <= 64'd1624553938728686361;
    6'd6: brom_out <= 64'd7147821265559899415;
    6'd7: brom_out <= 64'd3044098306375364542;
    6'd8: brom_out <= 64'd5976068779477487504;
    6'd9: brom_out <= 64'd3874323780530106533;
    6'd10: brom_out <= 64'd4066724171054462909;
    6'd11: brom_out <= 64'd2637886143940526168;
    6'd12: brom_out <= 64'd5792979130194094298;
    6'd13: brom_out <= 64'd2737158020017696281;
    6'd14: brom_out <= 64'd2803267708398697040;
    6'd15: brom_out <= 64'd1065160304167154726;
    6'd16: brom_out <= 64'd6551015095526749063;
    6'd17: brom_out <= 64'd8872444489401680815;
    6'd18: brom_out <= 64'd5908178380096272369;
    6'd19: brom_out <= 64'd3547627594494878621;
    6'd20: brom_out <= 64'd2991444385089030097;
    6'd21: brom_out <= 64'd9166670786663116443;
    6'd22: brom_out <= 64'd7646914504675205489;
    6'd23: brom_out <= 64'd4393262027419573708;
    6'd24: brom_out <= 64'd3392617565049336557;
    6'd25: brom_out <= 64'd5039744181953194803;
    6'd26: brom_out <= 64'd1002059954001900696;
    6'd27: brom_out <= 64'd9185509849420767578;
    6'd28: brom_out <= 64'd699101306064864663;
    6'd29: brom_out <= 64'd7923677684682802987;
    6'd30: brom_out <= 64'd1670791095363685175;
    6'd31: brom_out <= 64'd228503451388919711;
    default: brom_out <= 64'h1;
    endcase
end

generate
    if(DELAY == 1) begin
        assign b = brom_out;
    end
endgenerate

endmodule

//-------------------------------------------------------------------------------------------------

module tw_rom_6
#(
    parameter LOGN  = 6,
    parameter LOGQ  = 64,
    parameter DELAY = 1,
    parameter STAGE = 1
)(
    input            clk,
    input [LOGN-1:0] raddr,
    output[LOGQ-1:0] b
);

(* rom_style = "distributed" *)
reg [LOGQ-1:0] brom_out, brom_out2;

always @(posedge clk) begin
    case(raddr[STAGE-1:0])
    7'd0: brom_out <= 64'd9223372036854251519;
    7'd1: brom_out <= 64'd6984365454624050605;
    7'd2: brom_out <= 64'd8706294438413809553;
    7'd3: brom_out <= 64'd6158485483849164736;
    7'd4: brom_out <= 64'd5917339183240377480;
    7'd5: brom_out <= 64'd3950921523134993168;
    7'd6: brom_out <= 64'd4110363107264655732;
    7'd7: brom_out <= 64'd2194362728065833183;
    7'd8: brom_out <= 64'd2881966912403406253;
    7'd9: brom_out <= 64'd735439083491420630;
    7'd10: brom_out <= 64'd1624553938728686361;
    7'd11: brom_out <= 64'd5875474638474206446;
    7'd12: brom_out <= 64'd7147821265559899415;
    7'd13: brom_out <= 64'd8826561644056073004;
    7'd14: brom_out <= 64'd3044098306375364542;
    7'd15: brom_out <= 64'd3522401398456133729;
    7'd16: brom_out <= 64'd5976068779477487504;
    7'd17: brom_out <= 64'd8439932809411290039;
    7'd18: brom_out <= 64'd3874323780530106533;
    7'd19: brom_out <= 64'd1085106348447748099;
    7'd20: brom_out <= 64'd4066724171054462909;
    7'd21: brom_out <= 64'd8309796333647791448;
    7'd22: brom_out <= 64'd2637886143940526168;
    7'd23: brom_out <= 64'd4291000205908552613;
    7'd24: brom_out <= 64'd5792979130194094298;
    7'd25: brom_out <= 64'd5596038778869841895;
    7'd26: brom_out <= 64'd2737158020017696281;
    7'd27: brom_out <= 64'd6071971305117248446;
    7'd28: brom_out <= 64'd2803267708398697040;
    7'd29: brom_out <= 64'd3003943219615574075;
    7'd30: brom_out <= 64'd1065160304167154726;
    7'd31: brom_out <= 64'd4910995540748981844;
    7'd32: brom_out <= 64'd6551015095526749063;
    7'd33: brom_out <= 64'd284038871857826017;
    7'd34: brom_out <= 64'd8872444489401680815;
    7'd35: brom_out <= 64'd2669547459691193432;
    7'd36: brom_out <= 64'd5908178380096272369;
    7'd37: brom_out <= 64'd1687335542159875606;
    7'd38: brom_out <= 64'd3547627594494878621;
    7'd39: brom_out <= 64'd2468663283803736374;
    7'd40: brom_out <= 64'd2991444385089030097;
    7'd41: brom_out <= 64'd8124953238658307565;
    7'd42: brom_out <= 64'd9166670786663116443;
    7'd43: brom_out <= 64'd5654726277541044038;
    7'd44: brom_out <= 64'd7646914504675205489;
    7'd45: brom_out <= 64'd2141707773911427712;
    7'd46: brom_out <= 64'd4393262027419573708;
    7'd47: brom_out <= 64'd5729951333194461427;
    7'd48: brom_out <= 64'd3392617565049336557;
    7'd49: brom_out <= 64'd8216761589456164;
    7'd50: brom_out <= 64'd5039744181953194803;
    7'd51: brom_out <= 64'd1628906345678539120;
    7'd52: brom_out <= 64'd1002059954001900696;
    7'd53: brom_out <= 64'd4836003352449041316;
    7'd54: brom_out <= 64'd9185509849420767578;
    7'd55: brom_out <= 64'd9003279055065478956;
    7'd56: brom_out <= 64'd699101306064864663;
    7'd57: brom_out <= 64'd69843017785227084;
    7'd58: brom_out <= 64'd7923677684682802987;
    7'd59: brom_out <= 64'd5126845061066175356;
    7'd60: brom_out <= 64'd1670791095363685175;
    7'd61: brom_out <= 64'd8823464365455855293;
    7'd62: brom_out <= 64'd228503451388919711;
    7'd63: brom_out <= 64'd700730835196570872;
    default: brom_out <= 64'h1;
    endcase
end

generate
    if(DELAY == 1) begin
        assign b = brom_out;
    end
endgenerate

endmodule

//-------------------------------------------------------------------------------------------------

module tw_rom_7
#(
    parameter LOGN  = 7,
    parameter LOGQ  = 64,
    parameter DELAY = 1,
    parameter STAGE = 1
)(
    input            clk,
    input [LOGN-1:0] raddr,
    output[LOGQ-1:0] b
);

(* rom_style = "distributed" *)
reg [LOGQ-1:0] brom_out, brom_out2;

always @(posedge clk) begin
    case(raddr[STAGE-1:0])
    8'd0: brom_out <= 64'd9223372036854251519;
    8'd1: brom_out <= 64'd269998454485676360;
    8'd2: brom_out <= 64'd6984365454624050605;
    8'd3: brom_out <= 64'd5653377166457707394;
    8'd4: brom_out <= 64'd8706294438413809553;
    8'd5: brom_out <= 64'd6626061600160634657;
    8'd6: brom_out <= 64'd6158485483849164736;
    8'd7: brom_out <= 64'd7345482494331839697;
    8'd8: brom_out <= 64'd5917339183240377480;
    8'd9: brom_out <= 64'd8174323033676948403;
    8'd10: brom_out <= 64'd3950921523134993168;
    8'd11: brom_out <= 64'd4573453364429337213;
    8'd12: brom_out <= 64'd4110363107264655732;
    8'd13: brom_out <= 64'd8070303386396255336;
    8'd14: brom_out <= 64'd2194362728065833183;
    8'd15: brom_out <= 64'd6564530672913887453;
    8'd16: brom_out <= 64'd2881966912403406253;
    8'd17: brom_out <= 64'd1219064800028085468;
    8'd18: brom_out <= 64'd735439083491420630;
    8'd19: brom_out <= 64'd544940125055465581;
    8'd20: brom_out <= 64'd1624553938728686361;
    8'd21: brom_out <= 64'd2926075365041679386;
    8'd22: brom_out <= 64'd5875474638474206446;
    8'd23: brom_out <= 64'd6222003843073247882;
    8'd24: brom_out <= 64'd7147821265559899415;
    8'd25: brom_out <= 64'd4717392765204693644;
    8'd26: brom_out <= 64'd8826561644056073004;
    8'd27: brom_out <= 64'd3526492789053904424;
    8'd28: brom_out <= 64'd3044098306375364542;
    8'd29: brom_out <= 64'd221168427156668620;
    8'd30: brom_out <= 64'd3522401398456133729;
    8'd31: brom_out <= 64'd9025502593406216690;
    8'd32: brom_out <= 64'd5976068779477487504;
    8'd33: brom_out <= 64'd1271675644934090509;
    8'd34: brom_out <= 64'd8439932809411290039;
    8'd35: brom_out <= 64'd9036648888917473750;
    8'd36: brom_out <= 64'd3874323780530106533;
    8'd37: brom_out <= 64'd4363004334232094865;
    8'd38: brom_out <= 64'd1085106348447748099;
    8'd39: brom_out <= 64'd1403509903281381135;
    8'd40: brom_out <= 64'd4066724171054462909;
    8'd41: brom_out <= 64'd4710964611444245301;
    8'd42: brom_out <= 64'd8309796333647791448;
    8'd43: brom_out <= 64'd4441590473776765300;
    8'd44: brom_out <= 64'd2637886143940526168;
    8'd45: brom_out <= 64'd7086452204833135780;
    8'd46: brom_out <= 64'd4291000205908552613;
    8'd47: brom_out <= 64'd6665838607271236324;
    8'd48: brom_out <= 64'd5792979130194094298;
    8'd49: brom_out <= 64'd5318975219191802577;
    8'd50: brom_out <= 64'd5596038778869841895;
    8'd51: brom_out <= 64'd6458351418566661432;
    8'd52: brom_out <= 64'd2737158020017696281;
    8'd53: brom_out <= 64'd2216455649141208680;
    8'd54: brom_out <= 64'd6071971305117248446;
    8'd55: brom_out <= 64'd4050420130283138042;
    8'd56: brom_out <= 64'd2803267708398697040;
    8'd57: brom_out <= 64'd4083878445077305523;
    8'd58: brom_out <= 64'd3003943219615574075;
    8'd59: brom_out <= 64'd6019869478886392755;
    8'd60: brom_out <= 64'd1065160304167154726;
    8'd61: brom_out <= 64'd3598379093835291182;
    8'd62: brom_out <= 64'd4910995540748981844;
    8'd63: brom_out <= 64'd8856063189815385885;
    8'd64: brom_out <= 64'd6551015095526749063;
    8'd65: brom_out <= 64'd4040899244153570090;
    8'd66: brom_out <= 64'd284038871857826017;
    8'd67: brom_out <= 64'd2529239563039080875;
    8'd68: brom_out <= 64'd8872444489401680815;
    8'd69: brom_out <= 64'd2703826489472427745;
    8'd70: brom_out <= 64'd2669547459691193432;
    8'd71: brom_out <= 64'd538390155169630246;
    8'd72: brom_out <= 64'd5908178380096272369;
    8'd73: brom_out <= 64'd9076916340755116149;
    8'd74: brom_out <= 64'd1687335542159875606;
    8'd75: brom_out <= 64'd4938289008039594695;
    8'd76: brom_out <= 64'd3547627594494878621;
    8'd77: brom_out <= 64'd5944864576936445287;
    8'd78: brom_out <= 64'd2468663283803736374;
    8'd79: brom_out <= 64'd1178188298187125443;
    8'd80: brom_out <= 64'd2991444385089030097;
    8'd81: brom_out <= 64'd6281663284576107517;
    8'd82: brom_out <= 64'd8124953238658307565;
    8'd83: brom_out <= 64'd5782598045554155253;
    8'd84: brom_out <= 64'd9166670786663116443;
    8'd85: brom_out <= 64'd3115848091286679823;
    8'd86: brom_out <= 64'd5654726277541044038;
    8'd87: brom_out <= 64'd3558399091024426444;
    8'd88: brom_out <= 64'd7646914504675205489;
    8'd89: brom_out <= 64'd1555308162728177297;
    8'd90: brom_out <= 64'd2141707773911427712;
    8'd91: brom_out <= 64'd7010796944267998638;
    8'd92: brom_out <= 64'd4393262027419573708;
    8'd93: brom_out <= 64'd4919595983980879989;
    8'd94: brom_out <= 64'd5729951333194461427;
    8'd95: brom_out <= 64'd1376701315345052441;
    8'd96: brom_out <= 64'd3392617565049336557;
    8'd97: brom_out <= 64'd2263269548655216762;
    8'd98: brom_out <= 64'd8216761589456164;
    8'd99: brom_out <= 64'd8186964208105355814;
    8'd100: brom_out <= 64'd5039744181953194803;
    8'd101: brom_out <= 64'd5471972468712594632;
    8'd102: brom_out <= 64'd1628906345678539120;
    8'd103: brom_out <= 64'd3528090222809025860;
    8'd104: brom_out <= 64'd1002059954001900696;
    8'd105: brom_out <= 64'd307156682351195017;
    8'd106: brom_out <= 64'd4836003352449041316;
    8'd107: brom_out <= 64'd6436331060924184539;
    8'd108: brom_out <= 64'd9185509849420767578;
    8'd109: brom_out <= 64'd7995675456769788758;
    8'd110: brom_out <= 64'd9003279055065478956;
    8'd111: brom_out <= 64'd1827606411485443129;
    8'd112: brom_out <= 64'd699101306064864663;
    8'd113: brom_out <= 64'd5893272571222366297;
    8'd114: brom_out <= 64'd69843017785227084;
    8'd115: brom_out <= 64'd7645071031480098655;
    8'd116: brom_out <= 64'd7923677684682802987;
    8'd117: brom_out <= 64'd375356035198548383;
    8'd118: brom_out <= 64'd5126845061066175356;
    8'd119: brom_out <= 64'd796180145389681740;
    8'd120: brom_out <= 64'd1670791095363685175;
    8'd121: brom_out <= 64'd3280526131456603436;
    8'd122: brom_out <= 64'd8823464365455855293;
    8'd123: brom_out <= 64'd8323983203612776937;
    8'd124: brom_out <= 64'd228503451388919711;
    8'd125: brom_out <= 64'd7002130558985726630;
    8'd126: brom_out <= 64'd700730835196570872;
    8'd127: brom_out <= 64'd2113561489472542490;
    default: brom_out <= 64'h1;
    endcase
end

generate
    if(DELAY == 1) begin
        assign b = brom_out;
    end
endgenerate

endmodule

//-------------------------------------------------------------------------------------------------

module tw_rom_8
#(
    parameter LOGN  = 8,
    parameter LOGQ  = 64,
    parameter DELAY = 1,
    parameter STAGE = 1
)(
    input            clk,
    input [LOGN-1:0] raddr,
    output[LOGQ-1:0] b
);

(* ram_style = "block" *)
reg [LOGQ-1:0] brom_out, brom_out2;

always @(posedge clk) begin
    case(raddr[STAGE-1:0])
    9'd0: brom_out <= 64'd9223372036854251519;
    9'd1: brom_out <= 64'd1299456045732977605;
    9'd2: brom_out <= 64'd269998454485676360;
    9'd3: brom_out <= 64'd9033387621081412018;
    9'd4: brom_out <= 64'd6984365454624050605;
    9'd5: brom_out <= 64'd810060818546034655;
    9'd6: brom_out <= 64'd5653377166457707394;
    9'd7: brom_out <= 64'd8914698016797979130;
    9'd8: brom_out <= 64'd8706294438413809553;
    9'd9: brom_out <= 64'd1984480336129885140;
    9'd10: brom_out <= 64'd6626061600160634657;
    9'd11: brom_out <= 64'd6375267241083926885;
    9'd12: brom_out <= 64'd6158485483849164736;
    9'd13: brom_out <= 64'd2808688244394002011;
    9'd14: brom_out <= 64'd7345482494331839697;
    9'd15: brom_out <= 64'd8037037384829722617;
    9'd16: brom_out <= 64'd5917339183240377480;
    9'd17: brom_out <= 64'd3561119328844693546;
    9'd18: brom_out <= 64'd8174323033676948403;
    9'd19: brom_out <= 64'd2319035647868930894;
    9'd20: brom_out <= 64'd3950921523134993168;
    9'd21: brom_out <= 64'd3531419639158455240;
    9'd22: brom_out <= 64'd4573453364429337213;
    9'd23: brom_out <= 64'd3367056065757602806;
    9'd24: brom_out <= 64'd4110363107264655732;
    9'd25: brom_out <= 64'd5233426006749936404;
    9'd26: brom_out <= 64'd8070303386396255336;
    9'd27: brom_out <= 64'd5682374489572555945;
    9'd28: brom_out <= 64'd2194362728065833183;
    9'd29: brom_out <= 64'd240070673848085803;
    9'd30: brom_out <= 64'd6564530672913887453;
    9'd31: brom_out <= 64'd1907082839763808740;
    9'd32: brom_out <= 64'd2881966912403406253;
    9'd33: brom_out <= 64'd8852621130615879035;
    9'd34: brom_out <= 64'd1219064800028085468;
    9'd35: brom_out <= 64'd1865389637899575391;
    9'd36: brom_out <= 64'd735439083491420630;
    9'd37: brom_out <= 64'd4936662293846854616;
    9'd38: brom_out <= 64'd544940125055465581;
    9'd39: brom_out <= 64'd1845447672304840611;
    9'd40: brom_out <= 64'd1624553938728686361;
    9'd41: brom_out <= 64'd3586995478868233709;
    9'd42: brom_out <= 64'd2926075365041679386;
    9'd43: brom_out <= 64'd5712154480457087476;
    9'd44: brom_out <= 64'd5875474638474206446;
    9'd45: brom_out <= 64'd7289325041362829578;
    9'd46: brom_out <= 64'd6222003843073247882;
    9'd47: brom_out <= 64'd616529505270125954;
    9'd48: brom_out <= 64'd7147821265559899415;
    9'd49: brom_out <= 64'd3149227341269420724;
    9'd50: brom_out <= 64'd4717392765204693644;
    9'd51: brom_out <= 64'd4312120720500409507;
    9'd52: brom_out <= 64'd8826561644056073004;
    9'd53: brom_out <= 64'd7048641871031816;
    9'd54: brom_out <= 64'd3526492789053904424;
    9'd55: brom_out <= 64'd5311697839062869272;
    9'd56: brom_out <= 64'd3044098306375364542;
    9'd57: brom_out <= 64'd7940586545958498989;
    9'd58: brom_out <= 64'd221168427156668620;
    9'd59: brom_out <= 64'd5446263128435942946;
    9'd60: brom_out <= 64'd3522401398456133729;
    9'd61: brom_out <= 64'd7748187342122623094;
    9'd62: brom_out <= 64'd9025502593406216690;
    9'd63: brom_out <= 64'd4533570374417505243;
    9'd64: brom_out <= 64'd5976068779477487504;
    9'd65: brom_out <= 64'd593042282816257658;
    9'd66: brom_out <= 64'd1271675644934090509;
    9'd67: brom_out <= 64'd1177438167634269823;
    9'd68: brom_out <= 64'd8439932809411290039;
    9'd69: brom_out <= 64'd9170359323010223211;
    9'd70: brom_out <= 64'd9036648888917473750;
    9'd71: brom_out <= 64'd739218949392655402;
    9'd72: brom_out <= 64'd3874323780530106533;
    9'd73: brom_out <= 64'd5718867093180509803;
    9'd74: brom_out <= 64'd4363004334232094865;
    9'd75: brom_out <= 64'd7929071200947786101;
    9'd76: brom_out <= 64'd1085106348447748099;
    9'd77: brom_out <= 64'd809486194630696952;
    9'd78: brom_out <= 64'd1403509903281381135;
    9'd79: brom_out <= 64'd4619323584991910886;
    9'd80: brom_out <= 64'd4066724171054462909;
    9'd81: brom_out <= 64'd3603203538984367077;
    9'd82: brom_out <= 64'd4710964611444245301;
    9'd83: brom_out <= 64'd6828380608571071779;
    9'd84: brom_out <= 64'd8309796333647791448;
    9'd85: brom_out <= 64'd5684075750352032262;
    9'd86: brom_out <= 64'd4441590473776765300;
    9'd87: brom_out <= 64'd6707938413484059878;
    9'd88: brom_out <= 64'd2637886143940526168;
    9'd89: brom_out <= 64'd5320908759602881481;
    9'd90: brom_out <= 64'd7086452204833135780;
    9'd91: brom_out <= 64'd3372994486386929879;
    9'd92: brom_out <= 64'd4291000205908552613;
    9'd93: brom_out <= 64'd1232654478032123658;
    9'd94: brom_out <= 64'd6665838607271236324;
    9'd95: brom_out <= 64'd4070504440077246346;
    9'd96: brom_out <= 64'd5792979130194094298;
    9'd97: brom_out <= 64'd222968537858942369;
    9'd98: brom_out <= 64'd5318975219191802577;
    9'd99: brom_out <= 64'd5000944239179137954;
    9'd100: brom_out <= 64'd5596038778869841895;
    9'd101: brom_out <= 64'd3365288337767276247;
    9'd102: brom_out <= 64'd6458351418566661432;
    9'd103: brom_out <= 64'd5293457782313866956;
    9'd104: brom_out <= 64'd2737158020017696281;
    9'd105: brom_out <= 64'd5607163649712091882;
    9'd106: brom_out <= 64'd2216455649141208680;
    9'd107: brom_out <= 64'd1455837426791755297;
    9'd108: brom_out <= 64'd6071971305117248446;
    9'd109: brom_out <= 64'd2023644405886518221;
    9'd110: brom_out <= 64'd4050420130283138042;
    9'd111: brom_out <= 64'd5243772136807645099;
    9'd112: brom_out <= 64'd2803267708398697040;
    9'd113: brom_out <= 64'd1618067356643750162;
    9'd114: brom_out <= 64'd4083878445077305523;
    9'd115: brom_out <= 64'd7741923924364988008;
    9'd116: brom_out <= 64'd3003943219615574075;
    9'd117: brom_out <= 64'd2803062370827609981;
    9'd118: brom_out <= 64'd6019869478886392755;
    9'd119: brom_out <= 64'd5746142847633122703;
    9'd120: brom_out <= 64'd1065160304167154726;
    9'd121: brom_out <= 64'd8151167855892330172;
    9'd122: brom_out <= 64'd3598379093835291182;
    9'd123: brom_out <= 64'd4667723862850537194;
    9'd124: brom_out <= 64'd4910995540748981844;
    9'd125: brom_out <= 64'd9009408318896786413;
    9'd126: brom_out <= 64'd8856063189815385885;
    9'd127: brom_out <= 64'd4891968351182874667;
    9'd128: brom_out <= 64'd6551015095526749063;
    9'd129: brom_out <= 64'd3796382495133268725;
    9'd130: brom_out <= 64'd4040899244153570090;
    9'd131: brom_out <= 64'd5683041679221725246;
    9'd132: brom_out <= 64'd284038871857826017;
    9'd133: brom_out <= 64'd2554384204381077376;
    9'd134: brom_out <= 64'd2529239563039080875;
    9'd135: brom_out <= 64'd9106909176665937792;
    9'd136: brom_out <= 64'd8872444489401680815;
    9'd137: brom_out <= 64'd4613289516563687559;
    9'd138: brom_out <= 64'd2703826489472427745;
    9'd139: brom_out <= 64'd1952843272151728048;
    9'd140: brom_out <= 64'd2669547459691193432;
    9'd141: brom_out <= 64'd8345571030034495946;
    9'd142: brom_out <= 64'd538390155169630246;
    9'd143: brom_out <= 64'd4078971191093288272;
    9'd144: brom_out <= 64'd5908178380096272369;
    9'd145: brom_out <= 64'd4682857295746554344;
    9'd146: brom_out <= 64'd9076916340755116149;
    9'd147: brom_out <= 64'd5040843640203270416;
    9'd148: brom_out <= 64'd1687335542159875606;
    9'd149: brom_out <= 64'd8818463071528412136;
    9'd150: brom_out <= 64'd4938289008039594695;
    9'd151: brom_out <= 64'd6574977840107373503;
    9'd152: brom_out <= 64'd3547627594494878621;
    9'd153: brom_out <= 64'd57560180524151836;
    9'd154: brom_out <= 64'd5944864576936445287;
    9'd155: brom_out <= 64'd684639643803771175;
    9'd156: brom_out <= 64'd2468663283803736374;
    9'd157: brom_out <= 64'd1837680713908133646;
    9'd158: brom_out <= 64'd1178188298187125443;
    9'd159: brom_out <= 64'd5873106135293020355;
    9'd160: brom_out <= 64'd2991444385089030097;
    9'd161: brom_out <= 64'd1122397655549924356;
    9'd162: brom_out <= 64'd6281663284576107517;
    9'd163: brom_out <= 64'd8697599446790123293;
    9'd164: brom_out <= 64'd8124953238658307565;
    9'd165: brom_out <= 64'd4625294087119433729;
    9'd166: brom_out <= 64'd5782598045554155253;
    9'd167: brom_out <= 64'd5991059833680697521;
    9'd168: brom_out <= 64'd9166670786663116443;
    9'd169: brom_out <= 64'd7173654840489607776;
    9'd170: brom_out <= 64'd3115848091286679823;
    9'd171: brom_out <= 64'd750361034814781007;
    9'd172: brom_out <= 64'd5654726277541044038;
    9'd173: brom_out <= 64'd5208814341045079371;
    9'd174: brom_out <= 64'd3558399091024426444;
    9'd175: brom_out <= 64'd4764036910647300995;
    9'd176: brom_out <= 64'd7646914504675205489;
    9'd177: brom_out <= 64'd3065938557921374089;
    9'd178: brom_out <= 64'd1555308162728177297;
    9'd179: brom_out <= 64'd6550225160897858344;
    9'd180: brom_out <= 64'd2141707773911427712;
    9'd181: brom_out <= 64'd5418439566171715291;
    9'd182: brom_out <= 64'd7010796944267998638;
    9'd183: brom_out <= 64'd8692551628537520016;
    9'd184: brom_out <= 64'd4393262027419573708;
    9'd185: brom_out <= 64'd4159689793066360690;
    9'd186: brom_out <= 64'd4919595983980879989;
    9'd187: brom_out <= 64'd4919750730687193807;
    9'd188: brom_out <= 64'd5729951333194461427;
    9'd189: brom_out <= 64'd2240289491309476277;
    9'd190: brom_out <= 64'd1376701315345052441;
    9'd191: brom_out <= 64'd5939667306004532036;
    9'd192: brom_out <= 64'd3392617565049336557;
    9'd193: brom_out <= 64'd7479147464852913991;
    9'd194: brom_out <= 64'd2263269548655216762;
    9'd195: brom_out <= 64'd6982695801609760735;
    9'd196: brom_out <= 64'd8216761589456164;
    9'd197: brom_out <= 64'd6925371594294004533;
    9'd198: brom_out <= 64'd8186964208105355814;
    9'd199: brom_out <= 64'd6849437044168275747;
    9'd200: brom_out <= 64'd5039744181953194803;
    9'd201: brom_out <= 64'd3064309850488305304;
    9'd202: brom_out <= 64'd5471972468712594632;
    9'd203: brom_out <= 64'd6626178562688381462;
    9'd204: brom_out <= 64'd1628906345678539120;
    9'd205: brom_out <= 64'd7705829573832500897;
    9'd206: brom_out <= 64'd3528090222809025860;
    9'd207: brom_out <= 64'd8798316185508471405;
    9'd208: brom_out <= 64'd1002059954001900696;
    9'd209: brom_out <= 64'd1490887556607246244;
    9'd210: brom_out <= 64'd307156682351195017;
    9'd211: brom_out <= 64'd3107918471259441615;
    9'd212: brom_out <= 64'd4836003352449041316;
    9'd213: brom_out <= 64'd2923414615723271043;
    9'd214: brom_out <= 64'd6436331060924184539;
    9'd215: brom_out <= 64'd1641922973023157952;
    9'd216: brom_out <= 64'd9185509849420767578;
    9'd217: brom_out <= 64'd1546731779372361302;
    9'd218: brom_out <= 64'd7995675456769788758;
    9'd219: brom_out <= 64'd4849682055056439114;
    9'd220: brom_out <= 64'd9003279055065478956;
    9'd221: brom_out <= 64'd869826359180825983;
    9'd222: brom_out <= 64'd1827606411485443129;
    9'd223: brom_out <= 64'd7672998258368931866;
    9'd224: brom_out <= 64'd699101306064864663;
    9'd225: brom_out <= 64'd8219959792660589692;
    9'd226: brom_out <= 64'd5893272571222366297;
    9'd227: brom_out <= 64'd4439925312673350003;
    9'd228: brom_out <= 64'd69843017785227084;
    9'd229: brom_out <= 64'd8225172405297280263;
    9'd230: brom_out <= 64'd7645071031480098655;
    9'd231: brom_out <= 64'd5173422508798334624;
    9'd232: brom_out <= 64'd7923677684682802987;
    9'd233: brom_out <= 64'd2139689406997953411;
    9'd234: brom_out <= 64'd375356035198548383;
    9'd235: brom_out <= 64'd511527761999251354;
    9'd236: brom_out <= 64'd5126845061066175356;
    9'd237: brom_out <= 64'd9162350688835803463;
    9'd238: brom_out <= 64'd796180145389681740;
    9'd239: brom_out <= 64'd4119508171639317112;
    9'd240: brom_out <= 64'd1670791095363685175;
    9'd241: brom_out <= 64'd5989914729659460893;
    9'd242: brom_out <= 64'd3280526131456603436;
    9'd243: brom_out <= 64'd3615127351505505023;
    9'd244: brom_out <= 64'd8823464365455855293;
    9'd245: brom_out <= 64'd5003529372930301250;
    9'd246: brom_out <= 64'd8323983203612776937;
    9'd247: brom_out <= 64'd5423351720389833865;
    9'd248: brom_out <= 64'd228503451388919711;
    9'd249: brom_out <= 64'd498968785704607628;
    9'd250: brom_out <= 64'd7002130558985726630;
    9'd251: brom_out <= 64'd7471415495952780188;
    9'd252: brom_out <= 64'd700730835196570872;
    9'd253: brom_out <= 64'd8584995141337045279;
    9'd254: brom_out <= 64'd2113561489472542490;
    9'd255: brom_out <= 64'd7269045898348823146;
    default: brom_out <= 64'h1;
    endcase
end

generate
    if(DELAY == 1) begin
        assign b = brom_out;
    end
endgenerate

endmodule

//-------------------------------------------------------------------------------------------------

module tw_rom_9
#(
    parameter LOGN  = 9,
    parameter LOGQ  = 64,
    parameter DELAY = 1,
    parameter STAGE = 1
)(
    input            clk,
    input [LOGN-1:0] raddr,
    output[LOGQ-1:0] b
);

(* ram_style = "block" *)
reg [LOGQ-1:0] brom_out, brom_out2;

always @(posedge clk) begin
    case(raddr[STAGE-1:0])
    10'd0: brom_out <= 64'd9223372036854251519;
    10'd1: brom_out <= 64'd7605493872853681221;
    10'd2: brom_out <= 64'd1299456045732977605;
    10'd3: brom_out <= 64'd8213948439719346069;
    10'd4: brom_out <= 64'd269998454485676360;
    10'd5: brom_out <= 64'd7934371085285641861;
    10'd6: brom_out <= 64'd9033387621081412018;
    10'd7: brom_out <= 64'd4765886196678305331;
    10'd8: brom_out <= 64'd6984365454624050605;
    10'd9: brom_out <= 64'd2123066514724381883;
    10'd10: brom_out <= 64'd810060818546034655;
    10'd11: brom_out <= 64'd8581206737579399620;
    10'd12: brom_out <= 64'd5653377166457707394;
    10'd13: brom_out <= 64'd2299841007653134372;
    10'd14: brom_out <= 64'd8914698016797979130;
    10'd15: brom_out <= 64'd5779395201958353378;
    10'd16: brom_out <= 64'd8706294438413809553;
    10'd17: brom_out <= 64'd2509796222201502174;
    10'd18: brom_out <= 64'd1984480336129885140;
    10'd19: brom_out <= 64'd7152306933764292478;
    10'd20: brom_out <= 64'd6626061600160634657;
    10'd21: brom_out <= 64'd4332795524147639451;
    10'd22: brom_out <= 64'd6375267241083926885;
    10'd23: brom_out <= 64'd792297214988562254;
    10'd24: brom_out <= 64'd6158485483849164736;
    10'd25: brom_out <= 64'd1966154900029444318;
    10'd26: brom_out <= 64'd2808688244394002011;
    10'd27: brom_out <= 64'd7902540812321798218;
    10'd28: brom_out <= 64'd7345482494331839697;
    10'd29: brom_out <= 64'd299894953115934099;
    10'd30: brom_out <= 64'd8037037384829722617;
    10'd31: brom_out <= 64'd9104612624170912214;
    10'd32: brom_out <= 64'd5917339183240377480;
    10'd33: brom_out <= 64'd4392041727794040139;
    10'd34: brom_out <= 64'd3561119328844693546;
    10'd35: brom_out <= 64'd2908884142996516879;
    10'd36: brom_out <= 64'd8174323033676948403;
    10'd37: brom_out <= 64'd7153542761736184733;
    10'd38: brom_out <= 64'd2319035647868930894;
    10'd39: brom_out <= 64'd5900439431409958858;
    10'd40: brom_out <= 64'd3950921523134993168;
    10'd41: brom_out <= 64'd2162992210110465427;
    10'd42: brom_out <= 64'd3531419639158455240;
    10'd43: brom_out <= 64'd6297866057014224030;
    10'd44: brom_out <= 64'd4573453364429337213;
    10'd45: brom_out <= 64'd1287149587930120656;
    10'd46: brom_out <= 64'd3367056065757602806;
    10'd47: brom_out <= 64'd3883460632785907410;
    10'd48: brom_out <= 64'd4110363107264655732;
    10'd49: brom_out <= 64'd5549948750888088698;
    10'd50: brom_out <= 64'd5233426006749936404;
    10'd51: brom_out <= 64'd7125634071680409905;
    10'd52: brom_out <= 64'd8070303386396255336;
    10'd53: brom_out <= 64'd4346701462512900589;
    10'd54: brom_out <= 64'd5682374489572555945;
    10'd55: brom_out <= 64'd173114810237193158;
    10'd56: brom_out <= 64'd2194362728065833183;
    10'd57: brom_out <= 64'd401958369407258982;
    10'd58: brom_out <= 64'd240070673848085803;
    10'd59: brom_out <= 64'd1427846036265206780;
    10'd60: brom_out <= 64'd6564530672913887453;
    10'd61: brom_out <= 64'd3098083654159802861;
    10'd62: brom_out <= 64'd1907082839763808740;
    10'd63: brom_out <= 64'd3031844387819961827;
    10'd64: brom_out <= 64'd2881966912403406253;
    10'd65: brom_out <= 64'd2925409531261716840;
    10'd66: brom_out <= 64'd8852621130615879035;
    10'd67: brom_out <= 64'd270496797777326527;
    10'd68: brom_out <= 64'd1219064800028085468;
    10'd69: brom_out <= 64'd543577740076728061;
    10'd70: brom_out <= 64'd1865389637899575391;
    10'd71: brom_out <= 64'd7923340214113792441;
    10'd72: brom_out <= 64'd735439083491420630;
    10'd73: brom_out <= 64'd5356334136853441455;
    10'd74: brom_out <= 64'd4936662293846854616;
    10'd75: brom_out <= 64'd5689831925774807956;
    10'd76: brom_out <= 64'd544940125055465581;
    10'd77: brom_out <= 64'd1297536695137410486;
    10'd78: brom_out <= 64'd1845447672304840611;
    10'd79: brom_out <= 64'd2182902326656347159;
    10'd80: brom_out <= 64'd1624553938728686361;
    10'd81: brom_out <= 64'd3012117742719754636;
    10'd82: brom_out <= 64'd3586995478868233709;
    10'd83: brom_out <= 64'd2057313745147478637;
    10'd84: brom_out <= 64'd2926075365041679386;
    10'd85: brom_out <= 64'd7993764406966422987;
    10'd86: brom_out <= 64'd5712154480457087476;
    10'd87: brom_out <= 64'd3479065458090349436;
    10'd88: brom_out <= 64'd5875474638474206446;
    10'd89: brom_out <= 64'd6548403254923287631;
    10'd90: brom_out <= 64'd7289325041362829578;
    10'd91: brom_out <= 64'd1785088414017673288;
    10'd92: brom_out <= 64'd6222003843073247882;
    10'd93: brom_out <= 64'd1990992240235617717;
    10'd94: brom_out <= 64'd616529505270125954;
    10'd95: brom_out <= 64'd4535501105232824056;
    10'd96: brom_out <= 64'd7147821265559899415;
    10'd97: brom_out <= 64'd1598994064067110291;
    10'd98: brom_out <= 64'd3149227341269420724;
    10'd99: brom_out <= 64'd904660340594613265;
    10'd100: brom_out <= 64'd4717392765204693644;
    10'd101: brom_out <= 64'd4359339040815035935;
    10'd102: brom_out <= 64'd4312120720500409507;
    10'd103: brom_out <= 64'd749037117208255733;
    10'd104: brom_out <= 64'd8826561644056073004;
    10'd105: brom_out <= 64'd6153283181782085767;
    10'd106: brom_out <= 64'd7048641871031816;
    10'd107: brom_out <= 64'd3017602207931310620;
    10'd108: brom_out <= 64'd3526492789053904424;
    10'd109: brom_out <= 64'd489108130890476637;
    10'd110: brom_out <= 64'd5311697839062869272;
    10'd111: brom_out <= 64'd7009454947613216741;
    10'd112: brom_out <= 64'd3044098306375364542;
    10'd113: brom_out <= 64'd967392942188980461;
    10'd114: brom_out <= 64'd7940586545958498989;
    10'd115: brom_out <= 64'd8888883322669091370;
    10'd116: brom_out <= 64'd221168427156668620;
    10'd117: brom_out <= 64'd6954602674252549157;
    10'd118: brom_out <= 64'd5446263128435942946;
    10'd119: brom_out <= 64'd5301890443195662787;
    10'd120: brom_out <= 64'd3522401398456133729;
    10'd121: brom_out <= 64'd6985849834050000541;
    10'd122: brom_out <= 64'd7748187342122623094;
    10'd123: brom_out <= 64'd4187235956733982846;
    10'd124: brom_out <= 64'd9025502593406216690;
    10'd125: brom_out <= 64'd1744638522500329828;
    10'd126: brom_out <= 64'd4533570374417505243;
    10'd127: brom_out <= 64'd2914465977735506303;
    10'd128: brom_out <= 64'd5976068779477487504;
    10'd129: brom_out <= 64'd6061870125418198147;
    10'd130: brom_out <= 64'd593042282816257658;
    10'd131: brom_out <= 64'd5181330732459777477;
    10'd132: brom_out <= 64'd1271675644934090509;
    10'd133: brom_out <= 64'd8013822734360034103;
    10'd134: brom_out <= 64'd1177438167634269823;
    10'd135: brom_out <= 64'd6903674494547403458;
    10'd136: brom_out <= 64'd8439932809411290039;
    10'd137: brom_out <= 64'd8791519766434938211;
    10'd138: brom_out <= 64'd9170359323010223211;
    10'd139: brom_out <= 64'd4794628727443279888;
    10'd140: brom_out <= 64'd9036648888917473750;
    10'd141: brom_out <= 64'd994064848121607400;
    10'd142: brom_out <= 64'd739218949392655402;
    10'd143: brom_out <= 64'd7256022154194582960;
    10'd144: brom_out <= 64'd3874323780530106533;
    10'd145: brom_out <= 64'd6928014622416298408;
    10'd146: brom_out <= 64'd5718867093180509803;
    10'd147: brom_out <= 64'd8433488676012520446;
    10'd148: brom_out <= 64'd4363004334232094865;
    10'd149: brom_out <= 64'd1021589499332145736;
    10'd150: brom_out <= 64'd7929071200947786101;
    10'd151: brom_out <= 64'd2663302601066611311;
    10'd152: brom_out <= 64'd1085106348447748099;
    10'd153: brom_out <= 64'd853076967703601242;
    10'd154: brom_out <= 64'd809486194630696952;
    10'd155: brom_out <= 64'd6179534021270744021;
    10'd156: brom_out <= 64'd1403509903281381135;
    10'd157: brom_out <= 64'd3510417462984237944;
    10'd158: brom_out <= 64'd4619323584991910886;
    10'd159: brom_out <= 64'd6415125647473131768;
    10'd160: brom_out <= 64'd4066724171054462909;
    10'd161: brom_out <= 64'd1611893969776626643;
    10'd162: brom_out <= 64'd3603203538984367077;
    10'd163: brom_out <= 64'd8041554051968754776;
    10'd164: brom_out <= 64'd4710964611444245301;
    10'd165: brom_out <= 64'd3118801396391702857;
    10'd166: brom_out <= 64'd6828380608571071779;
    10'd167: brom_out <= 64'd8127637090793435339;
    10'd168: brom_out <= 64'd8309796333647791448;
    10'd169: brom_out <= 64'd7940540358792163042;
    10'd170: brom_out <= 64'd5684075750352032262;
    10'd171: brom_out <= 64'd6468256505106281226;
    10'd172: brom_out <= 64'd4441590473776765300;
    10'd173: brom_out <= 64'd8634381596625442610;
    10'd174: brom_out <= 64'd6707938413484059878;
    10'd175: brom_out <= 64'd8077069361822515059;
    10'd176: brom_out <= 64'd2637886143940526168;
    10'd177: brom_out <= 64'd4132551802894357262;
    10'd178: brom_out <= 64'd5320908759602881481;
    10'd179: brom_out <= 64'd6222808144614635014;
    10'd180: brom_out <= 64'd7086452204833135780;
    10'd181: brom_out <= 64'd5695358218414993869;
    10'd182: brom_out <= 64'd3372994486386929879;
    10'd183: brom_out <= 64'd3022260544642597516;
    10'd184: brom_out <= 64'd4291000205908552613;
    10'd185: brom_out <= 64'd7819977419197775899;
    10'd186: brom_out <= 64'd1232654478032123658;
    10'd187: brom_out <= 64'd7099443897569798910;
    10'd188: brom_out <= 64'd6665838607271236324;
    10'd189: brom_out <= 64'd1297339388260599077;
    10'd190: brom_out <= 64'd4070504440077246346;
    10'd191: brom_out <= 64'd7603550242876584926;
    10'd192: brom_out <= 64'd5792979130194094298;
    10'd193: brom_out <= 64'd4452291514428477137;
    10'd194: brom_out <= 64'd222968537858942369;
    10'd195: brom_out <= 64'd6650157038584548422;
    10'd196: brom_out <= 64'd5318975219191802577;
    10'd197: brom_out <= 64'd4110541742333500737;
    10'd198: brom_out <= 64'd5000944239179137954;
    10'd199: brom_out <= 64'd1059548844895002697;
    10'd200: brom_out <= 64'd5596038778869841895;
    10'd201: brom_out <= 64'd7803653637595225642;
    10'd202: brom_out <= 64'd3365288337767276247;
    10'd203: brom_out <= 64'd5892854050328892876;
    10'd204: brom_out <= 64'd6458351418566661432;
    10'd205: brom_out <= 64'd4456208975303951299;
    10'd206: brom_out <= 64'd5293457782313866956;
    10'd207: brom_out <= 64'd2351375173829121150;
    10'd208: brom_out <= 64'd2737158020017696281;
    10'd209: brom_out <= 64'd2487979883454043411;
    10'd210: brom_out <= 64'd5607163649712091882;
    10'd211: brom_out <= 64'd6229174968075775630;
    10'd212: brom_out <= 64'd2216455649141208680;
    10'd213: brom_out <= 64'd1314986123610772272;
    10'd214: brom_out <= 64'd1455837426791755297;
    10'd215: brom_out <= 64'd1701272341948035267;
    10'd216: brom_out <= 64'd6071971305117248446;
    10'd217: brom_out <= 64'd8108747189882628079;
    10'd218: brom_out <= 64'd2023644405886518221;
    10'd219: brom_out <= 64'd6396414439770314375;
    10'd220: brom_out <= 64'd4050420130283138042;
    10'd221: brom_out <= 64'd7977797132770592727;
    10'd222: brom_out <= 64'd5243772136807645099;
    10'd223: brom_out <= 64'd2314914454150418602;
    10'd224: brom_out <= 64'd2803267708398697040;
    10'd225: brom_out <= 64'd8376944661285632772;
    10'd226: brom_out <= 64'd1618067356643750162;
    10'd227: brom_out <= 64'd2784388700362841711;
    10'd228: brom_out <= 64'd4083878445077305523;
    10'd229: brom_out <= 64'd6337223876791081151;
    10'd230: brom_out <= 64'd7741923924364988008;
    10'd231: brom_out <= 64'd2215604315896092670;
    10'd232: brom_out <= 64'd3003943219615574075;
    10'd233: brom_out <= 64'd1382872280811698552;
    10'd234: brom_out <= 64'd2803062370827609981;
    10'd235: brom_out <= 64'd7700372050315114363;
    10'd236: brom_out <= 64'd6019869478886392755;
    10'd237: brom_out <= 64'd6761610796267635122;
    10'd238: brom_out <= 64'd5746142847633122703;
    10'd239: brom_out <= 64'd3130462232530454679;
    10'd240: brom_out <= 64'd1065160304167154726;
    10'd241: brom_out <= 64'd6953881865491377297;
    10'd242: brom_out <= 64'd8151167855892330172;
    10'd243: brom_out <= 64'd4976637449741390052;
    10'd244: brom_out <= 64'd3598379093835291182;
    10'd245: brom_out <= 64'd3659981058207187100;
    10'd246: brom_out <= 64'd4667723862850537194;
    10'd247: brom_out <= 64'd9119962653750090131;
    10'd248: brom_out <= 64'd4910995540748981844;
    10'd249: brom_out <= 64'd6432548891759686389;
    10'd250: brom_out <= 64'd9009408318896786413;
    10'd251: brom_out <= 64'd5184317378868141180;
    10'd252: brom_out <= 64'd8856063189815385885;
    10'd253: brom_out <= 64'd5590202575696230393;
    10'd254: brom_out <= 64'd4891968351182874667;
    10'd255: brom_out <= 64'd5145477708918912727;
    10'd256: brom_out <= 64'd6551015095526749063;
    10'd257: brom_out <= 64'd8652315721870189437;
    10'd258: brom_out <= 64'd3796382495133268725;
    10'd259: brom_out <= 64'd15243861875148476;
    10'd260: brom_out <= 64'd4040899244153570090;
    10'd261: brom_out <= 64'd2240211916433264831;
    10'd262: brom_out <= 64'd5683041679221725246;
    10'd263: brom_out <= 64'd8708624953667028585;
    10'd264: brom_out <= 64'd284038871857826017;
    10'd265: brom_out <= 64'd7096948766236504610;
    10'd266: brom_out <= 64'd2554384204381077376;
    10'd267: brom_out <= 64'd6463166748036722757;
    10'd268: brom_out <= 64'd2529239563039080875;
    10'd269: brom_out <= 64'd3847574256498121621;
    10'd270: brom_out <= 64'd9106909176665937792;
    10'd271: brom_out <= 64'd111332146913263916;
    10'd272: brom_out <= 64'd8872444489401680815;
    10'd273: brom_out <= 64'd2343344652186686753;
    10'd274: brom_out <= 64'd4613289516563687559;
    10'd275: brom_out <= 64'd6832924728641330482;
    10'd276: brom_out <= 64'd2703826489472427745;
    10'd277: brom_out <= 64'd3227682425404315158;
    10'd278: brom_out <= 64'd1952843272151728048;
    10'd279: brom_out <= 64'd7104270022735541970;
    10'd280: brom_out <= 64'd2669547459691193432;
    10'd281: brom_out <= 64'd4585039786213636068;
    10'd282: brom_out <= 64'd8345571030034495946;
    10'd283: brom_out <= 64'd6017550373169230213;
    10'd284: brom_out <= 64'd538390155169630246;
    10'd285: brom_out <= 64'd1458993785378647509;
    10'd286: brom_out <= 64'd4078971191093288272;
    10'd287: brom_out <= 64'd4583234557640069978;
    10'd288: brom_out <= 64'd5908178380096272369;
    10'd289: brom_out <= 64'd7993813175591520204;
    10'd290: brom_out <= 64'd4682857295746554344;
    10'd291: brom_out <= 64'd8934879803166669689;
    10'd292: brom_out <= 64'd9076916340755116149;
    10'd293: brom_out <= 64'd5024898852976039286;
    10'd294: brom_out <= 64'd5040843640203270416;
    10'd295: brom_out <= 64'd4506204908127599502;
    10'd296: brom_out <= 64'd1687335542159875606;
    10'd297: brom_out <= 64'd6854317339658753350;
    10'd298: brom_out <= 64'd8818463071528412136;
    10'd299: brom_out <= 64'd7284478466022368184;
    10'd300: brom_out <= 64'd4938289008039594695;
    10'd301: brom_out <= 64'd3688954750038363726;
    10'd302: brom_out <= 64'd6574977840107373503;
    10'd303: brom_out <= 64'd821107918729627811;
    10'd304: brom_out <= 64'd3547627594494878621;
    10'd305: brom_out <= 64'd1549287551893278911;
    10'd306: brom_out <= 64'd57560180524151836;
    10'd307: brom_out <= 64'd7831437647304356508;
    10'd308: brom_out <= 64'd5944864576936445287;
    10'd309: brom_out <= 64'd5078991997579173257;
    10'd310: brom_out <= 64'd684639643803771175;
    10'd311: brom_out <= 64'd3340259218302706899;
    10'd312: brom_out <= 64'd2468663283803736374;
    10'd313: brom_out <= 64'd5798824876843371582;
    10'd314: brom_out <= 64'd1837680713908133646;
    10'd315: brom_out <= 64'd2036591841189774695;
    10'd316: brom_out <= 64'd1178188298187125443;
    10'd317: brom_out <= 64'd3110559949174149380;
    10'd318: brom_out <= 64'd5873106135293020355;
    10'd319: brom_out <= 64'd8803778985884906727;
    10'd320: brom_out <= 64'd2991444385089030097;
    10'd321: brom_out <= 64'd4183299227927339195;
    10'd322: brom_out <= 64'd1122397655549924356;
    10'd323: brom_out <= 64'd2527297775950676908;
    10'd324: brom_out <= 64'd6281663284576107517;
    10'd325: brom_out <= 64'd7533491753178725717;
    10'd326: brom_out <= 64'd8697599446790123293;
    10'd327: brom_out <= 64'd235142833563334451;
    10'd328: brom_out <= 64'd8124953238658307565;
    10'd329: brom_out <= 64'd5808776274764837854;
    10'd330: brom_out <= 64'd4625294087119433729;
    10'd331: brom_out <= 64'd75966845172534173;
    10'd332: brom_out <= 64'd5782598045554155253;
    10'd333: brom_out <= 64'd7870108581299121483;
    10'd334: brom_out <= 64'd5991059833680697521;
    10'd335: brom_out <= 64'd8100294372597586432;
    10'd336: brom_out <= 64'd9166670786663116443;
    10'd337: brom_out <= 64'd7083423175763586691;
    10'd338: brom_out <= 64'd7173654840489607776;
    10'd339: brom_out <= 64'd1947243181919420491;
    10'd340: brom_out <= 64'd3115848091286679823;
    10'd341: brom_out <= 64'd5226535173943436928;
    10'd342: brom_out <= 64'd750361034814781007;
    10'd343: brom_out <= 64'd3592198641247208794;
    10'd344: brom_out <= 64'd5654726277541044038;
    10'd345: brom_out <= 64'd4510264232516592952;
    10'd346: brom_out <= 64'd5208814341045079371;
    10'd347: brom_out <= 64'd5551115908770807940;
    10'd348: brom_out <= 64'd3558399091024426444;
    10'd349: brom_out <= 64'd1491544262489362891;
    10'd350: brom_out <= 64'd4764036910647300995;
    10'd351: brom_out <= 64'd9197868711120196895;
    10'd352: brom_out <= 64'd7646914504675205489;
    10'd353: brom_out <= 64'd5713577346046003020;
    10'd354: brom_out <= 64'd3065938557921374089;
    10'd355: brom_out <= 64'd2744296939060575530;
    10'd356: brom_out <= 64'd1555308162728177297;
    10'd357: brom_out <= 64'd220088159844794260;
    10'd358: brom_out <= 64'd6550225160897858344;
    10'd359: brom_out <= 64'd5490294517849368108;
    10'd360: brom_out <= 64'd2141707773911427712;
    10'd361: brom_out <= 64'd7593220218804307867;
    10'd362: brom_out <= 64'd5418439566171715291;
    10'd363: brom_out <= 64'd4249431574386262900;
    10'd364: brom_out <= 64'd7010796944267998638;
    10'd365: brom_out <= 64'd7135696680823117604;
    10'd366: brom_out <= 64'd8692551628537520016;
    10'd367: brom_out <= 64'd4824069180043442917;
    10'd368: brom_out <= 64'd4393262027419573708;
    10'd369: brom_out <= 64'd8893614490103508778;
    10'd370: brom_out <= 64'd4159689793066360690;
    10'd371: brom_out <= 64'd654752926994167022;
    10'd372: brom_out <= 64'd4919595983980879989;
    10'd373: brom_out <= 64'd2816403948006974041;
    10'd374: brom_out <= 64'd4919750730687193807;
    10'd375: brom_out <= 64'd4413826527383477878;
    10'd376: brom_out <= 64'd5729951333194461427;
    10'd377: brom_out <= 64'd8743332571195579934;
    10'd378: brom_out <= 64'd2240289491309476277;
    10'd379: brom_out <= 64'd2173356542276770935;
    10'd380: brom_out <= 64'd1376701315345052441;
    10'd381: brom_out <= 64'd3167756150689666531;
    10'd382: brom_out <= 64'd5939667306004532036;
    10'd383: brom_out <= 64'd2935114005611711057;
    10'd384: brom_out <= 64'd3392617565049336557;
    10'd385: brom_out <= 64'd2230049327513614869;
    10'd386: brom_out <= 64'd7479147464852913991;
    10'd387: brom_out <= 64'd7538107808473199530;
    10'd388: brom_out <= 64'd2263269548655216762;
    10'd389: brom_out <= 64'd6798664954031634633;
    10'd390: brom_out <= 64'd6982695801609760735;
    10'd391: brom_out <= 64'd6068442745462420874;
    10'd392: brom_out <= 64'd8216761589456164;
    10'd393: brom_out <= 64'd9102413699342598757;
    10'd394: brom_out <= 64'd6925371594294004533;
    10'd395: brom_out <= 64'd1568136098664689522;
    10'd396: brom_out <= 64'd8186964208105355814;
    10'd397: brom_out <= 64'd1676869911627098617;
    10'd398: brom_out <= 64'd6849437044168275747;
    10'd399: brom_out <= 64'd8444867741212273661;
    10'd400: brom_out <= 64'd5039744181953194803;
    10'd401: brom_out <= 64'd3468732936118861906;
    10'd402: brom_out <= 64'd3064309850488305304;
    10'd403: brom_out <= 64'd391518006782257654;
    10'd404: brom_out <= 64'd5471972468712594632;
    10'd405: brom_out <= 64'd8395167631823199941;
    10'd406: brom_out <= 64'd6626178562688381462;
    10'd407: brom_out <= 64'd9209536114756024834;
    10'd408: brom_out <= 64'd1628906345678539120;
    10'd409: brom_out <= 64'd4368700210148671551;
    10'd410: brom_out <= 64'd7705829573832500897;
    10'd411: brom_out <= 64'd4934228471949137670;
    10'd412: brom_out <= 64'd3528090222809025860;
    10'd413: brom_out <= 64'd1258669831230654444;
    10'd414: brom_out <= 64'd8798316185508471405;
    10'd415: brom_out <= 64'd6154077313509807261;
    10'd416: brom_out <= 64'd1002059954001900696;
    10'd417: brom_out <= 64'd2757773614559033666;
    10'd418: brom_out <= 64'd1490887556607246244;
    10'd419: brom_out <= 64'd7104811893195087792;
    10'd420: brom_out <= 64'd307156682351195017;
    10'd421: brom_out <= 64'd8730278730941939396;
    10'd422: brom_out <= 64'd3107918471259441615;
    10'd423: brom_out <= 64'd6460685242337216620;
    10'd424: brom_out <= 64'd4836003352449041316;
    10'd425: brom_out <= 64'd8051296741047110195;
    10'd426: brom_out <= 64'd2923414615723271043;
    10'd427: brom_out <= 64'd8026629062288902533;
    10'd428: brom_out <= 64'd6436331060924184539;
    10'd429: brom_out <= 64'd6733707155866364304;
    10'd430: brom_out <= 64'd1641922973023157952;
    10'd431: brom_out <= 64'd4681773058202772675;
    10'd432: brom_out <= 64'd9185509849420767578;
    10'd433: brom_out <= 64'd6230952056441481807;
    10'd434: brom_out <= 64'd1546731779372361302;
    10'd435: brom_out <= 64'd1790792280522562723;
    10'd436: brom_out <= 64'd7995675456769788758;
    10'd437: brom_out <= 64'd198235807530720187;
    10'd438: brom_out <= 64'd4849682055056439114;
    10'd439: brom_out <= 64'd9160052455972965925;
    10'd440: brom_out <= 64'd9003279055065478956;
    10'd441: brom_out <= 64'd5011986474190685475;
    10'd442: brom_out <= 64'd869826359180825983;
    10'd443: brom_out <= 64'd6630229277550940928;
    10'd444: brom_out <= 64'd1827606411485443129;
    10'd445: brom_out <= 64'd6949147395764538964;
    10'd446: brom_out <= 64'd7672998258368931866;
    10'd447: brom_out <= 64'd7530731249570041776;
    10'd448: brom_out <= 64'd699101306064864663;
    10'd449: brom_out <= 64'd655123889431899961;
    10'd450: brom_out <= 64'd8219959792660589692;
    10'd451: brom_out <= 64'd8543830174923091154;
    10'd452: brom_out <= 64'd5893272571222366297;
    10'd453: brom_out <= 64'd2015889517693822068;
    10'd454: brom_out <= 64'd4439925312673350003;
    10'd455: brom_out <= 64'd4798734633597747276;
    10'd456: brom_out <= 64'd69843017785227084;
    10'd457: brom_out <= 64'd8247980103556855667;
    10'd458: brom_out <= 64'd8225172405297280263;
    10'd459: brom_out <= 64'd976868090527140556;
    10'd460: brom_out <= 64'd7645071031480098655;
    10'd461: brom_out <= 64'd5140288024937627165;
    10'd462: brom_out <= 64'd5173422508798334624;
    10'd463: brom_out <= 64'd2600298912569494844;
    10'd464: brom_out <= 64'd7923677684682802987;
    10'd465: brom_out <= 64'd2275953281661646751;
    10'd466: brom_out <= 64'd2139689406997953411;
    10'd467: brom_out <= 64'd3729764982569583119;
    10'd468: brom_out <= 64'd375356035198548383;
    10'd469: brom_out <= 64'd4961919869715327681;
    10'd470: brom_out <= 64'd511527761999251354;
    10'd471: brom_out <= 64'd5412893724914022449;
    10'd472: brom_out <= 64'd5126845061066175356;
    10'd473: brom_out <= 64'd6181066534637459237;
    10'd474: brom_out <= 64'd9162350688835803463;
    10'd475: brom_out <= 64'd841949363898762459;
    10'd476: brom_out <= 64'd796180145389681740;
    10'd477: brom_out <= 64'd6881112568257936145;
    10'd478: brom_out <= 64'd4119508171639317112;
    10'd479: brom_out <= 64'd4523573697502160143;
    10'd480: brom_out <= 64'd1670791095363685175;
    10'd481: brom_out <= 64'd6268445540391799960;
    10'd482: brom_out <= 64'd5989914729659460893;
    10'd483: brom_out <= 64'd8498706274306490892;
    10'd484: brom_out <= 64'd3280526131456603436;
    10'd485: brom_out <= 64'd881381962624186811;
    10'd486: brom_out <= 64'd3615127351505505023;
    10'd487: brom_out <= 64'd6148609810148795929;
    10'd488: brom_out <= 64'd8823464365455855293;
    10'd489: brom_out <= 64'd5139097896322553033;
    10'd490: brom_out <= 64'd5003529372930301250;
    10'd491: brom_out <= 64'd3363566323249637328;
    10'd492: brom_out <= 64'd8323983203612776937;
    10'd493: brom_out <= 64'd3740576396473059045;
    10'd494: brom_out <= 64'd5423351720389833865;
    10'd495: brom_out <= 64'd5408302969401217960;
    10'd496: brom_out <= 64'd228503451388919711;
    10'd497: brom_out <= 64'd6913883903315781469;
    10'd498: brom_out <= 64'd498968785704607628;
    10'd499: brom_out <= 64'd3083280881619226755;
    10'd500: brom_out <= 64'd7002130558985726630;
    10'd501: brom_out <= 64'd3016980039216328962;
    10'd502: brom_out <= 64'd7471415495952780188;
    10'd503: brom_out <= 64'd9117660520541870682;
    10'd504: brom_out <= 64'd700730835196570872;
    10'd505: brom_out <= 64'd7087203385146507098;
    10'd506: brom_out <= 64'd8584995141337045279;
    10'd507: brom_out <= 64'd6918964554399920495;
    10'd508: brom_out <= 64'd2113561489472542490;
    10'd509: brom_out <= 64'd3835383961103183096;
    10'd510: brom_out <= 64'd7269045898348823146;
    10'd511: brom_out <= 64'd8634110784643349010;
    default: brom_out <= 64'h1;
    endcase
end

generate
    if(DELAY == 1) begin
        assign b = brom_out;
    end
endgenerate

endmodule

//-------------------------------------------------------------------------------------------------

module tw_rom_10
#(
    parameter LOGN  = 10,
    parameter LOGQ  = 64,
    parameter DELAY = 1,
    parameter STAGE = 1
)(
    input            clk,
    input [LOGN-1:0] raddr,
    output[LOGQ-1:0] b
);

(* ram_style = "block" *)
reg [LOGQ-1:0] brom_out, brom_out2;

always @(posedge clk) begin
    case(raddr[STAGE-1:0])
    11'd0: brom_out <= 64'd9223372036854251519;
    11'd1: brom_out <= 64'd6012871302989280084;
    11'd2: brom_out <= 64'd7605493872853681221;
    11'd3: brom_out <= 64'd3127052517479868225;
    11'd4: brom_out <= 64'd1299456045732977605;
    11'd5: brom_out <= 64'd9150256334426485369;
    11'd6: brom_out <= 64'd8213948439719346069;
    11'd7: brom_out <= 64'd6825597430088558793;
    11'd8: brom_out <= 64'd269998454485676360;
    11'd9: brom_out <= 64'd2564423744727517704;
    11'd10: brom_out <= 64'd7934371085285641861;
    11'd11: brom_out <= 64'd7153207102067290344;
    11'd12: brom_out <= 64'd9033387621081412018;
    11'd13: brom_out <= 64'd3293074636399430213;
    11'd14: brom_out <= 64'd4765886196678305331;
    11'd15: brom_out <= 64'd5112583091541522973;
    11'd16: brom_out <= 64'd6984365454624050605;
    11'd17: brom_out <= 64'd2273617654662494576;
    11'd18: brom_out <= 64'd2123066514724381883;
    11'd19: brom_out <= 64'd2567313654253520317;
    11'd20: brom_out <= 64'd810060818546034655;
    11'd21: brom_out <= 64'd6588969549873072984;
    11'd22: brom_out <= 64'd8581206737579399620;
    11'd23: brom_out <= 64'd7820318430984191122;
    11'd24: brom_out <= 64'd5653377166457707394;
    11'd25: brom_out <= 64'd2934009396408142147;
    11'd26: brom_out <= 64'd2299841007653134372;
    11'd27: brom_out <= 64'd1287674294028378649;
    11'd28: brom_out <= 64'd8914698016797979130;
    11'd29: brom_out <= 64'd4290018412507268451;
    11'd30: brom_out <= 64'd5779395201958353378;
    11'd31: brom_out <= 64'd8710174058585331351;
    11'd32: brom_out <= 64'd8706294438413809553;
    11'd33: brom_out <= 64'd6756792246403704650;
    11'd34: brom_out <= 64'd2509796222201502174;
    11'd35: brom_out <= 64'd1467033842096743702;
    11'd36: brom_out <= 64'd1984480336129885140;
    11'd37: brom_out <= 64'd5411415188401616703;
    11'd38: brom_out <= 64'd7152306933764292478;
    11'd39: brom_out <= 64'd8367416970837404480;
    11'd40: brom_out <= 64'd6626061600160634657;
    11'd41: brom_out <= 64'd1408687539684857079;
    11'd42: brom_out <= 64'd4332795524147639451;
    11'd43: brom_out <= 64'd6891504871357446422;
    11'd44: brom_out <= 64'd6375267241083926885;
    11'd45: brom_out <= 64'd7586867602903602858;
    11'd46: brom_out <= 64'd792297214988562254;
    11'd47: brom_out <= 64'd7058677087284092182;
    11'd48: brom_out <= 64'd6158485483849164736;
    11'd49: brom_out <= 64'd5266916899250488660;
    11'd50: brom_out <= 64'd1966154900029444318;
    11'd51: brom_out <= 64'd1215003878949612048;
    11'd52: brom_out <= 64'd2808688244394002011;
    11'd53: brom_out <= 64'd3851039626226392450;
    11'd54: brom_out <= 64'd7902540812321798218;
    11'd55: brom_out <= 64'd6004430279489338680;
    11'd56: brom_out <= 64'd7345482494331839697;
    11'd57: brom_out <= 64'd4218632253198916038;
    11'd58: brom_out <= 64'd299894953115934099;
    11'd59: brom_out <= 64'd1821424608084578998;
    11'd60: brom_out <= 64'd8037037384829722617;
    11'd61: brom_out <= 64'd4110036900460384796;
    11'd62: brom_out <= 64'd9104612624170912214;
    11'd63: brom_out <= 64'd1547693224024900634;
    11'd64: brom_out <= 64'd5917339183240377480;
    11'd65: brom_out <= 64'd8498480881154740865;
    11'd66: brom_out <= 64'd4392041727794040139;
    11'd67: brom_out <= 64'd6475240946856553091;
    11'd68: brom_out <= 64'd3561119328844693546;
    11'd69: brom_out <= 64'd5569609541362591627;
    11'd70: brom_out <= 64'd2908884142996516879;
    11'd71: brom_out <= 64'd3495906847793555496;
    11'd72: brom_out <= 64'd8174323033676948403;
    11'd73: brom_out <= 64'd8346874721972884401;
    11'd74: brom_out <= 64'd7153542761736184733;
    11'd75: brom_out <= 64'd9036614214691043214;
    11'd76: brom_out <= 64'd2319035647868930894;
    11'd77: brom_out <= 64'd1331680507007219705;
    11'd78: brom_out <= 64'd5900439431409958858;
    11'd79: brom_out <= 64'd8944063972887106670;
    11'd80: brom_out <= 64'd3950921523134993168;
    11'd81: brom_out <= 64'd2884516234218684811;
    11'd82: brom_out <= 64'd2162992210110465427;
    11'd83: brom_out <= 64'd7920402332462387511;
    11'd84: brom_out <= 64'd3531419639158455240;
    11'd85: brom_out <= 64'd7396774219033937672;
    11'd86: brom_out <= 64'd6297866057014224030;
    11'd87: brom_out <= 64'd1188483528343374386;
    11'd88: brom_out <= 64'd4573453364429337213;
    11'd89: brom_out <= 64'd6252329300465472480;
    11'd90: brom_out <= 64'd1287149587930120656;
    11'd91: brom_out <= 64'd5698207036020272794;
    11'd92: brom_out <= 64'd3367056065757602806;
    11'd93: brom_out <= 64'd118243567567768095;
    11'd94: brom_out <= 64'd3883460632785907410;
    11'd95: brom_out <= 64'd4486934250525894693;
    11'd96: brom_out <= 64'd4110363107264655732;
    11'd97: brom_out <= 64'd4514892859148397044;
    11'd98: brom_out <= 64'd5549948750888088698;
    11'd99: brom_out <= 64'd2943321537520600659;
    11'd100: brom_out <= 64'd5233426006749936404;
    11'd101: brom_out <= 64'd5747717726212286166;
    11'd102: brom_out <= 64'd7125634071680409905;
    11'd103: brom_out <= 64'd4614122134803297477;
    11'd104: brom_out <= 64'd8070303386396255336;
    11'd105: brom_out <= 64'd8117367890929318445;
    11'd106: brom_out <= 64'd4346701462512900589;
    11'd107: brom_out <= 64'd7783606212229745263;
    11'd108: brom_out <= 64'd5682374489572555945;
    11'd109: brom_out <= 64'd880050980480071141;
    11'd110: brom_out <= 64'd173114810237193158;
    11'd111: brom_out <= 64'd5314247580215590840;
    11'd112: brom_out <= 64'd2194362728065833183;
    11'd113: brom_out <= 64'd7403262497201993765;
    11'd114: brom_out <= 64'd401958369407258982;
    11'd115: brom_out <= 64'd4151717614504932492;
    11'd116: brom_out <= 64'd240070673848085803;
    11'd117: brom_out <= 64'd4057166001169818856;
    11'd118: brom_out <= 64'd1427846036265206780;
    11'd119: brom_out <= 64'd5295131112655049137;
    11'd120: brom_out <= 64'd6564530672913887453;
    11'd121: brom_out <= 64'd3866632472152804465;
    11'd122: brom_out <= 64'd3098083654159802861;
    11'd123: brom_out <= 64'd3063481684957609078;
    11'd124: brom_out <= 64'd1907082839763808740;
    11'd125: brom_out <= 64'd1468430662791236228;
    11'd126: brom_out <= 64'd3031844387819961827;
    11'd127: brom_out <= 64'd1396316958451531348;
    11'd128: brom_out <= 64'd2881966912403406253;
    11'd129: brom_out <= 64'd9146187461299601623;
    11'd130: brom_out <= 64'd2925409531261716840;
    11'd131: brom_out <= 64'd4304180803912282259;
    11'd132: brom_out <= 64'd8852621130615879035;
    11'd133: brom_out <= 64'd4848840577486999766;
    11'd134: brom_out <= 64'd270496797777326527;
    11'd135: brom_out <= 64'd6083010805285052716;
    11'd136: brom_out <= 64'd1219064800028085468;
    11'd137: brom_out <= 64'd6306667576969932326;
    11'd138: brom_out <= 64'd543577740076728061;
    11'd139: brom_out <= 64'd4091222591604623441;
    11'd140: brom_out <= 64'd1865389637899575391;
    11'd141: brom_out <= 64'd2862891865227566885;
    11'd142: brom_out <= 64'd7923340214113792441;
    11'd143: brom_out <= 64'd4822434129781452362;
    11'd144: brom_out <= 64'd735439083491420630;
    11'd145: brom_out <= 64'd8701208384429075876;
    11'd146: brom_out <= 64'd5356334136853441455;
    11'd147: brom_out <= 64'd2004505146951275140;
    11'd148: brom_out <= 64'd4936662293846854616;
    11'd149: brom_out <= 64'd695669619354178199;
    11'd150: brom_out <= 64'd5689831925774807956;
    11'd151: brom_out <= 64'd1189038338221773258;
    11'd152: brom_out <= 64'd544940125055465581;
    11'd153: brom_out <= 64'd2331992164875830888;
    11'd154: brom_out <= 64'd1297536695137410486;
    11'd155: brom_out <= 64'd4174433604295068968;
    11'd156: brom_out <= 64'd1845447672304840611;
    11'd157: brom_out <= 64'd7530083780768442237;
    11'd158: brom_out <= 64'd2182902326656347159;
    11'd159: brom_out <= 64'd7697402264257745017;
    11'd160: brom_out <= 64'd1624553938728686361;
    11'd161: brom_out <= 64'd2235543617824736075;
    11'd162: brom_out <= 64'd3012117742719754636;
    11'd163: brom_out <= 64'd8395034085139528506;
    11'd164: brom_out <= 64'd3586995478868233709;
    11'd165: brom_out <= 64'd5121098992128955161;
    11'd166: brom_out <= 64'd2057313745147478637;
    11'd167: brom_out <= 64'd5160625525529957528;
    11'd168: brom_out <= 64'd2926075365041679386;
    11'd169: brom_out <= 64'd3516066647433260551;
    11'd170: brom_out <= 64'd7993764406966422987;
    11'd171: brom_out <= 64'd8037258735659770483;
    11'd172: brom_out <= 64'd5712154480457087476;
    11'd173: brom_out <= 64'd3018928514936204385;
    11'd174: brom_out <= 64'd3479065458090349436;
    11'd175: brom_out <= 64'd1585371721068583241;
    11'd176: brom_out <= 64'd5875474638474206446;
    11'd177: brom_out <= 64'd4515128673629883118;
    11'd178: brom_out <= 64'd6548403254923287631;
    11'd179: brom_out <= 64'd4752592209480917425;
    11'd180: brom_out <= 64'd7289325041362829578;
    11'd181: brom_out <= 64'd6185725345812273456;
    11'd182: brom_out <= 64'd1785088414017673288;
    11'd183: brom_out <= 64'd4798463378767722612;
    11'd184: brom_out <= 64'd6222003843073247882;
    11'd185: brom_out <= 64'd3324417521285869935;
    11'd186: brom_out <= 64'd1990992240235617717;
    11'd187: brom_out <= 64'd8528027318223251457;
    11'd188: brom_out <= 64'd616529505270125954;
    11'd189: brom_out <= 64'd1960716502804548672;
    11'd190: brom_out <= 64'd4535501105232824056;
    11'd191: brom_out <= 64'd2293080637268173952;
    11'd192: brom_out <= 64'd7147821265559899415;
    11'd193: brom_out <= 64'd8249092968287330570;
    11'd194: brom_out <= 64'd1598994064067110291;
    11'd195: brom_out <= 64'd6446311831687328438;
    11'd196: brom_out <= 64'd3149227341269420724;
    11'd197: brom_out <= 64'd2519301650103661960;
    11'd198: brom_out <= 64'd904660340594613265;
    11'd199: brom_out <= 64'd3412151563337741352;
    11'd200: brom_out <= 64'd4717392765204693644;
    11'd201: brom_out <= 64'd865268308687100412;
    11'd202: brom_out <= 64'd4359339040815035935;
    11'd203: brom_out <= 64'd5458238346969861276;
    11'd204: brom_out <= 64'd4312120720500409507;
    11'd205: brom_out <= 64'd3241756220799506222;
    11'd206: brom_out <= 64'd749037117208255733;
    11'd207: brom_out <= 64'd8021309328199436730;
    11'd208: brom_out <= 64'd8826561644056073004;
    11'd209: brom_out <= 64'd6492936536869808625;
    11'd210: brom_out <= 64'd6153283181782085767;
    11'd211: brom_out <= 64'd3042490808619695370;
    11'd212: brom_out <= 64'd7048641871031816;
    11'd213: brom_out <= 64'd6938251047297990533;
    11'd214: brom_out <= 64'd3017602207931310620;
    11'd215: brom_out <= 64'd6526255316566008010;
    11'd216: brom_out <= 64'd3526492789053904424;
    11'd217: brom_out <= 64'd1097341705165972594;
    11'd218: brom_out <= 64'd489108130890476637;
    11'd219: brom_out <= 64'd9168100354083393324;
    11'd220: brom_out <= 64'd5311697839062869272;
    11'd221: brom_out <= 64'd3754010688254048597;
    11'd222: brom_out <= 64'd7009454947613216741;
    11'd223: brom_out <= 64'd1722163249877292090;
    11'd224: brom_out <= 64'd3044098306375364542;
    11'd225: brom_out <= 64'd3652792854953481228;
    11'd226: brom_out <= 64'd967392942188980461;
    11'd227: brom_out <= 64'd494499881005363032;
    11'd228: brom_out <= 64'd7940586545958498989;
    11'd229: brom_out <= 64'd5108575401283476645;
    11'd230: brom_out <= 64'd8888883322669091370;
    11'd231: brom_out <= 64'd2151578802008365031;
    11'd232: brom_out <= 64'd221168427156668620;
    11'd233: brom_out <= 64'd7985210005529564458;
    11'd234: brom_out <= 64'd6954602674252549157;
    11'd235: brom_out <= 64'd3877069780779427166;
    11'd236: brom_out <= 64'd5446263128435942946;
    11'd237: brom_out <= 64'd8162841956676165738;
    11'd238: brom_out <= 64'd5301890443195662787;
    11'd239: brom_out <= 64'd1123132456013002459;
    11'd240: brom_out <= 64'd3522401398456133729;
    11'd241: brom_out <= 64'd4785516395754103712;
    11'd242: brom_out <= 64'd6985849834050000541;
    11'd243: brom_out <= 64'd6520183508896026597;
    11'd244: brom_out <= 64'd7748187342122623094;
    11'd245: brom_out <= 64'd6590112200699224071;
    11'd246: brom_out <= 64'd4187235956733982846;
    11'd247: brom_out <= 64'd4635191165656492150;
    11'd248: brom_out <= 64'd9025502593406216690;
    11'd249: brom_out <= 64'd5775523390321313615;
    11'd250: brom_out <= 64'd1744638522500329828;
    11'd251: brom_out <= 64'd3651945852037892795;
    11'd252: brom_out <= 64'd4533570374417505243;
    11'd253: brom_out <= 64'd9097630694651455464;
    11'd254: brom_out <= 64'd2914465977735506303;
    11'd255: brom_out <= 64'd8074623464407446434;
    11'd256: brom_out <= 64'd5976068779477487504;
    11'd257: brom_out <= 64'd6744020006969895307;
    11'd258: brom_out <= 64'd6061870125418198147;
    11'd259: brom_out <= 64'd8927943298820454076;
    11'd260: brom_out <= 64'd593042282816257658;
    11'd261: brom_out <= 64'd2799537887104471251;
    11'd262: brom_out <= 64'd5181330732459777477;
    11'd263: brom_out <= 64'd2187018093810691720;
    11'd264: brom_out <= 64'd1271675644934090509;
    11'd265: brom_out <= 64'd8522993162440537939;
    11'd266: brom_out <= 64'd8013822734360034103;
    11'd267: brom_out <= 64'd5541375517500192895;
    11'd268: brom_out <= 64'd1177438167634269823;
    11'd269: brom_out <= 64'd7698250944354989161;
    11'd270: brom_out <= 64'd6903674494547403458;
    11'd271: brom_out <= 64'd5401614836719703272;
    11'd272: brom_out <= 64'd8439932809411290039;
    11'd273: brom_out <= 64'd5152644225124011089;
    11'd274: brom_out <= 64'd8791519766434938211;
    11'd275: brom_out <= 64'd2868266086180312958;
    11'd276: brom_out <= 64'd9170359323010223211;
    11'd277: brom_out <= 64'd4765782474432323605;
    11'd278: brom_out <= 64'd4794628727443279888;
    11'd279: brom_out <= 64'd4633112736508198766;
    11'd280: brom_out <= 64'd9036648888917473750;
    11'd281: brom_out <= 64'd8336322066205089657;
    11'd282: brom_out <= 64'd994064848121607400;
    11'd283: brom_out <= 64'd5410674334166473286;
    11'd284: brom_out <= 64'd739218949392655402;
    11'd285: brom_out <= 64'd8105253848644364450;
    11'd286: brom_out <= 64'd7256022154194582960;
    11'd287: brom_out <= 64'd2464563482745670645;
    11'd288: brom_out <= 64'd3874323780530106533;
    11'd289: brom_out <= 64'd6351756831470743006;
    11'd290: brom_out <= 64'd6928014622416298408;
    11'd291: brom_out <= 64'd7747822092528642924;
    11'd292: brom_out <= 64'd5718867093180509803;
    11'd293: brom_out <= 64'd8252964877799973406;
    11'd294: brom_out <= 64'd8433488676012520446;
    11'd295: brom_out <= 64'd1481999355516963175;
    11'd296: brom_out <= 64'd4363004334232094865;
    11'd297: brom_out <= 64'd7137177962332868154;
    11'd298: brom_out <= 64'd1021589499332145736;
    11'd299: brom_out <= 64'd2857441601682776678;
    11'd300: brom_out <= 64'd7929071200947786101;
    11'd301: brom_out <= 64'd2703396381905810774;
    11'd302: brom_out <= 64'd2663302601066611311;
    11'd303: brom_out <= 64'd6034460869506398985;
    11'd304: brom_out <= 64'd1085106348447748099;
    11'd305: brom_out <= 64'd7280577718007746774;
    11'd306: brom_out <= 64'd853076967703601242;
    11'd307: brom_out <= 64'd8765870513679473211;
    11'd308: brom_out <= 64'd809486194630696952;
    11'd309: brom_out <= 64'd6768544696756439421;
    11'd310: brom_out <= 64'd6179534021270744021;
    11'd311: brom_out <= 64'd8658919390669651664;
    11'd312: brom_out <= 64'd1403509903281381135;
    11'd313: brom_out <= 64'd4551293125869120088;
    11'd314: brom_out <= 64'd3510417462984237944;
    11'd315: brom_out <= 64'd7524025148374291789;
    11'd316: brom_out <= 64'd4619323584991910886;
    11'd317: brom_out <= 64'd6326125611953081505;
    11'd318: brom_out <= 64'd6415125647473131768;
    11'd319: brom_out <= 64'd6658739335726264481;
    11'd320: brom_out <= 64'd4066724171054462909;
    11'd321: brom_out <= 64'd548261701981485419;
    11'd322: brom_out <= 64'd1611893969776626643;
    11'd323: brom_out <= 64'd9004572314107590138;
    11'd324: brom_out <= 64'd3603203538984367077;
    11'd325: brom_out <= 64'd2805030511231525764;
    11'd326: brom_out <= 64'd8041554051968754776;
    11'd327: brom_out <= 64'd4806777613109574958;
    11'd328: brom_out <= 64'd4710964611444245301;
    11'd329: brom_out <= 64'd6926030477489072308;
    11'd330: brom_out <= 64'd3118801396391702857;
    11'd331: brom_out <= 64'd6265810223453665551;
    11'd332: brom_out <= 64'd6828380608571071779;
    11'd333: brom_out <= 64'd1512800906605612428;
    11'd334: brom_out <= 64'd8127637090793435339;
    11'd335: brom_out <= 64'd4414284518212157732;
    11'd336: brom_out <= 64'd8309796333647791448;
    11'd337: brom_out <= 64'd6457789071063052555;
    11'd338: brom_out <= 64'd7940540358792163042;
    11'd339: brom_out <= 64'd3823809497424801247;
    11'd340: brom_out <= 64'd5684075750352032262;
    11'd341: brom_out <= 64'd1415882188212200225;
    11'd342: brom_out <= 64'd6468256505106281226;
    11'd343: brom_out <= 64'd5300966512209250050;
    11'd344: brom_out <= 64'd4441590473776765300;
    11'd345: brom_out <= 64'd787340924847783803;
    11'd346: brom_out <= 64'd8634381596625442610;
    11'd347: brom_out <= 64'd7704688953664041795;
    11'd348: brom_out <= 64'd6707938413484059878;
    11'd349: brom_out <= 64'd1689924925158498949;
    11'd350: brom_out <= 64'd8077069361822515059;
    11'd351: brom_out <= 64'd6919778738676338510;
    11'd352: brom_out <= 64'd2637886143940526168;
    11'd353: brom_out <= 64'd7047875822701595031;
    11'd354: brom_out <= 64'd4132551802894357262;
    11'd355: brom_out <= 64'd7687396513344217400;
    11'd356: brom_out <= 64'd5320908759602881481;
    11'd357: brom_out <= 64'd8135317976049821842;
    11'd358: brom_out <= 64'd6222808144614635014;
    11'd359: brom_out <= 64'd5991839321352371775;
    11'd360: brom_out <= 64'd7086452204833135780;
    11'd361: brom_out <= 64'd1213734665504106333;
    11'd362: brom_out <= 64'd5695358218414993869;
    11'd363: brom_out <= 64'd8240076708661524496;
    11'd364: brom_out <= 64'd3372994486386929879;
    11'd365: brom_out <= 64'd4519341334859734073;
    11'd366: brom_out <= 64'd3022260544642597516;
    11'd367: brom_out <= 64'd6353718731862795407;
    11'd368: brom_out <= 64'd4291000205908552613;
    11'd369: brom_out <= 64'd7224435870105783327;
    11'd370: brom_out <= 64'd7819977419197775899;
    11'd371: brom_out <= 64'd7149484177775971227;
    11'd372: brom_out <= 64'd1232654478032123658;
    11'd373: brom_out <= 64'd196307236251518595;
    11'd374: brom_out <= 64'd7099443897569798910;
    11'd375: brom_out <= 64'd1364531386125093388;
    11'd376: brom_out <= 64'd6665838607271236324;
    11'd377: brom_out <= 64'd3633365094721677201;
    11'd378: brom_out <= 64'd1297339388260599077;
    11'd379: brom_out <= 64'd4041634879120597886;
    11'd380: brom_out <= 64'd4070504440077246346;
    11'd381: brom_out <= 64'd5917399405983790504;
    11'd382: brom_out <= 64'd7603550242876584926;
    11'd383: brom_out <= 64'd7094683365482870580;
    11'd384: brom_out <= 64'd5792979130194094298;
    11'd385: brom_out <= 64'd1390063910113207289;
    11'd386: brom_out <= 64'd4452291514428477137;
    11'd387: brom_out <= 64'd7817367043308214467;
    11'd388: brom_out <= 64'd222968537858942369;
    11'd389: brom_out <= 64'd1539629244627310107;
    11'd390: brom_out <= 64'd6650157038584548422;
    11'd391: brom_out <= 64'd2456301622261705551;
    11'd392: brom_out <= 64'd5318975219191802577;
    11'd393: brom_out <= 64'd8995741913985100290;
    11'd394: brom_out <= 64'd4110541742333500737;
    11'd395: brom_out <= 64'd7055503816228831091;
    11'd396: brom_out <= 64'd5000944239179137954;
    11'd397: brom_out <= 64'd5215707159989682948;
    11'd398: brom_out <= 64'd1059548844895002697;
    11'd399: brom_out <= 64'd5359119263554810248;
    11'd400: brom_out <= 64'd5596038778869841895;
    11'd401: brom_out <= 64'd1852954710699492504;
    11'd402: brom_out <= 64'd7803653637595225642;
    11'd403: brom_out <= 64'd4446551631123665655;
    11'd404: brom_out <= 64'd3365288337767276247;
    11'd405: brom_out <= 64'd6519885780090122409;
    11'd406: brom_out <= 64'd5892854050328892876;
    11'd407: brom_out <= 64'd2086211756656440867;
    11'd408: brom_out <= 64'd6458351418566661432;
    11'd409: brom_out <= 64'd2721341105491390085;
    11'd410: brom_out <= 64'd4456208975303951299;
    11'd411: brom_out <= 64'd5852786553912777685;
    11'd412: brom_out <= 64'd5293457782313866956;
    11'd413: brom_out <= 64'd1503390632805335282;
    11'd414: brom_out <= 64'd2351375173829121150;
    11'd415: brom_out <= 64'd8759164961417563512;
    11'd416: brom_out <= 64'd2737158020017696281;
    11'd417: brom_out <= 64'd6640287097552321424;
    11'd418: brom_out <= 64'd2487979883454043411;
    11'd419: brom_out <= 64'd17521832455993642;
    11'd420: brom_out <= 64'd5607163649712091882;
    11'd421: brom_out <= 64'd4217348036314092382;
    11'd422: brom_out <= 64'd6229174968075775630;
    11'd423: brom_out <= 64'd2051998054788366270;
    11'd424: brom_out <= 64'd2216455649141208680;
    11'd425: brom_out <= 64'd6796227057672368420;
    11'd426: brom_out <= 64'd1314986123610772272;
    11'd427: brom_out <= 64'd5880920423784685274;
    11'd428: brom_out <= 64'd1455837426791755297;
    11'd429: brom_out <= 64'd6481798364871042424;
    11'd430: brom_out <= 64'd1701272341948035267;
    11'd431: brom_out <= 64'd1168596851321766456;
    11'd432: brom_out <= 64'd6071971305117248446;
    11'd433: brom_out <= 64'd211205323560102598;
    11'd434: brom_out <= 64'd8108747189882628079;
    11'd435: brom_out <= 64'd962867634407305569;
    11'd436: brom_out <= 64'd2023644405886518221;
    11'd437: brom_out <= 64'd8948912045682648319;
    11'd438: brom_out <= 64'd6396414439770314375;
    11'd439: brom_out <= 64'd6259526245218962991;
    11'd440: brom_out <= 64'd4050420130283138042;
    11'd441: brom_out <= 64'd6160499120912117934;
    11'd442: brom_out <= 64'd7977797132770592727;
    11'd443: brom_out <= 64'd6552355050471698204;
    11'd444: brom_out <= 64'd5243772136807645099;
    11'd445: brom_out <= 64'd3651142297411659187;
    11'd446: brom_out <= 64'd2314914454150418602;
    11'd447: brom_out <= 64'd801305510105442737;
    11'd448: brom_out <= 64'd2803267708398697040;
    11'd449: brom_out <= 64'd4568079005623157455;
    11'd450: brom_out <= 64'd8376944661285632772;
    11'd451: brom_out <= 64'd8566281893646113;
    11'd452: brom_out <= 64'd1618067356643750162;
    11'd453: brom_out <= 64'd3507173358449499779;
    11'd454: brom_out <= 64'd2784388700362841711;
    11'd455: brom_out <= 64'd6295273620685999449;
    11'd456: brom_out <= 64'd4083878445077305523;
    11'd457: brom_out <= 64'd2848313604941519881;
    11'd458: brom_out <= 64'd6337223876791081151;
    11'd459: brom_out <= 64'd7990560214861353583;
    11'd460: brom_out <= 64'd7741923924364988008;
    11'd461: brom_out <= 64'd1144176920185415535;
    11'd462: brom_out <= 64'd2215604315896092670;
    11'd463: brom_out <= 64'd2608525535082964773;
    11'd464: brom_out <= 64'd3003943219615574075;
    11'd465: brom_out <= 64'd47740789800497965;
    11'd466: brom_out <= 64'd1382872280811698552;
    11'd467: brom_out <= 64'd1901574174662490027;
    11'd468: brom_out <= 64'd2803062370827609981;
    11'd469: brom_out <= 64'd1992283337758212979;
    11'd470: brom_out <= 64'd7700372050315114363;
    11'd471: brom_out <= 64'd2875223919672073068;
    11'd472: brom_out <= 64'd6019869478886392755;
    11'd473: brom_out <= 64'd7140722186488696864;
    11'd474: brom_out <= 64'd6761610796267635122;
    11'd475: brom_out <= 64'd3287964157657373940;
    11'd476: brom_out <= 64'd5746142847633122703;
    11'd477: brom_out <= 64'd3343459330700479572;
    11'd478: brom_out <= 64'd3130462232530454679;
    11'd479: brom_out <= 64'd6889879677402930206;
    11'd480: brom_out <= 64'd1065160304167154726;
    11'd481: brom_out <= 64'd8625960684678229166;
    11'd482: brom_out <= 64'd6953881865491377297;
    11'd483: brom_out <= 64'd1707361404853655714;
    11'd484: brom_out <= 64'd8151167855892330172;
    11'd485: brom_out <= 64'd4633933436842356737;
    11'd486: brom_out <= 64'd4976637449741390052;
    11'd487: brom_out <= 64'd6447223936141958870;
    11'd488: brom_out <= 64'd3598379093835291182;
    11'd489: brom_out <= 64'd3473787664538686576;
    11'd490: brom_out <= 64'd3659981058207187100;
    11'd491: brom_out <= 64'd8632467951852587989;
    11'd492: brom_out <= 64'd4667723862850537194;
    11'd493: brom_out <= 64'd3936667969893923919;
    11'd494: brom_out <= 64'd9119962653750090131;
    11'd495: brom_out <= 64'd168302224660410828;
    11'd496: brom_out <= 64'd4910995540748981844;
    11'd497: brom_out <= 64'd3657039766247532725;
    11'd498: brom_out <= 64'd6432548891759686389;
    11'd499: brom_out <= 64'd9123574294358671657;
    11'd500: brom_out <= 64'd9009408318896786413;
    11'd501: brom_out <= 64'd3633265221550976288;
    11'd502: brom_out <= 64'd5184317378868141180;
    11'd503: brom_out <= 64'd6244689180377020923;
    11'd504: brom_out <= 64'd8856063189815385885;
    11'd505: brom_out <= 64'd1118592617708714057;
    11'd506: brom_out <= 64'd5590202575696230393;
    11'd507: brom_out <= 64'd3794573246885287845;
    11'd508: brom_out <= 64'd4891968351182874667;
    11'd509: brom_out <= 64'd8063678981840380015;
    11'd510: brom_out <= 64'd5145477708918912727;
    11'd511: brom_out <= 64'd7920910159561005345;
    11'd512: brom_out <= 64'd6551015095526749063;
    11'd513: brom_out <= 64'd8288530531944855590;
    11'd514: brom_out <= 64'd8652315721870189437;
    11'd515: brom_out <= 64'd6914660438246835908;
    11'd516: brom_out <= 64'd3796382495133268725;
    11'd517: brom_out <= 64'd2726913976235435110;
    11'd518: brom_out <= 64'd15243861875148476;
    11'd519: brom_out <= 64'd4148280298264435145;
    11'd520: brom_out <= 64'd4040899244153570090;
    11'd521: brom_out <= 64'd4512365403662406081;
    11'd522: brom_out <= 64'd2240211916433264831;
    11'd523: brom_out <= 64'd7160540774931803866;
    11'd524: brom_out <= 64'd5683041679221725246;
    11'd525: brom_out <= 64'd9206702681534441482;
    11'd526: brom_out <= 64'd8708624953667028585;
    11'd527: brom_out <= 64'd7835211644950567469;
    11'd528: brom_out <= 64'd284038871857826017;
    11'd529: brom_out <= 64'd1445608483214028307;
    11'd530: brom_out <= 64'd7096948766236504610;
    11'd531: brom_out <= 64'd1778468342386166084;
    11'd532: brom_out <= 64'd2554384204381077376;
    11'd533: brom_out <= 64'd7537176118984402773;
    11'd534: brom_out <= 64'd6463166748036722757;
    11'd535: brom_out <= 64'd7664280676247221904;
    11'd536: brom_out <= 64'd2529239563039080875;
    11'd537: brom_out <= 64'd5407047594096528025;
    11'd538: brom_out <= 64'd3847574256498121621;
    11'd539: brom_out <= 64'd8373705960209865750;
    11'd540: brom_out <= 64'd9106909176665937792;
    11'd541: brom_out <= 64'd1100339483998246003;
    11'd542: brom_out <= 64'd111332146913263916;
    11'd543: brom_out <= 64'd849306692269551679;
    11'd544: brom_out <= 64'd8872444489401680815;
    11'd545: brom_out <= 64'd6943865764417683064;
    11'd546: brom_out <= 64'd2343344652186686753;
    11'd547: brom_out <= 64'd4751890286330071625;
    11'd548: brom_out <= 64'd4613289516563687559;
    11'd549: brom_out <= 64'd806771516604876704;
    11'd550: brom_out <= 64'd6832924728641330482;
    11'd551: brom_out <= 64'd6060747830154195747;
    11'd552: brom_out <= 64'd2703826489472427745;
    11'd553: brom_out <= 64'd3163609927867779470;
    11'd554: brom_out <= 64'd3227682425404315158;
    11'd555: brom_out <= 64'd5069629123053312106;
    11'd556: brom_out <= 64'd1952843272151728048;
    11'd557: brom_out <= 64'd5757481406149589238;
    11'd558: brom_out <= 64'd7104270022735541970;
    11'd559: brom_out <= 64'd812235029203875617;
    11'd560: brom_out <= 64'd2669547459691193432;
    11'd561: brom_out <= 64'd1709606027938467824;
    11'd562: brom_out <= 64'd4585039786213636068;
    11'd563: brom_out <= 64'd5269356158780504864;
    11'd564: brom_out <= 64'd8345571030034495946;
    11'd565: brom_out <= 64'd5711684474143641757;
    11'd566: brom_out <= 64'd6017550373169230213;
    11'd567: brom_out <= 64'd8871767897380268353;
    11'd568: brom_out <= 64'd538390155169630246;
    11'd569: brom_out <= 64'd7452519829483945138;
    11'd570: brom_out <= 64'd1458993785378647509;
    11'd571: brom_out <= 64'd6524722060171723622;
    11'd572: brom_out <= 64'd4078971191093288272;
    11'd573: brom_out <= 64'd6501664496823873080;
    11'd574: brom_out <= 64'd4583234557640069978;
    11'd575: brom_out <= 64'd6382089802135409144;
    11'd576: brom_out <= 64'd5908178380096272369;
    11'd577: brom_out <= 64'd9103463721653978408;
    11'd578: brom_out <= 64'd7993813175591520204;
    11'd579: brom_out <= 64'd3032208211650146388;
    11'd580: brom_out <= 64'd4682857295746554344;
    11'd581: brom_out <= 64'd3139435852145256442;
    11'd582: brom_out <= 64'd8934879803166669689;
    11'd583: brom_out <= 64'd6846824846681755777;
    11'd584: brom_out <= 64'd9076916340755116149;
    11'd585: brom_out <= 64'd6610810496821611972;
    11'd586: brom_out <= 64'd5024898852976039286;
    11'd587: brom_out <= 64'd5041872014433074100;
    11'd588: brom_out <= 64'd5040843640203270416;
    11'd589: brom_out <= 64'd789422816571225780;
    11'd590: brom_out <= 64'd4506204908127599502;
    11'd591: brom_out <= 64'd4822808530417619233;
    11'd592: brom_out <= 64'd1687335542159875606;
    11'd593: brom_out <= 64'd9135823465542849361;
    11'd594: brom_out <= 64'd6854317339658753350;
    11'd595: brom_out <= 64'd7125835522680848670;
    11'd596: brom_out <= 64'd8818463071528412136;
    11'd597: brom_out <= 64'd5992435799082823388;
    11'd598: brom_out <= 64'd7284478466022368184;
    11'd599: brom_out <= 64'd176563187302484685;
    11'd600: brom_out <= 64'd4938289008039594695;
    11'd601: brom_out <= 64'd5802647509516054700;
    11'd602: brom_out <= 64'd3688954750038363726;
    11'd603: brom_out <= 64'd287090937624021185;
    11'd604: brom_out <= 64'd6574977840107373503;
    11'd605: brom_out <= 64'd7077564256689660660;
    11'd606: brom_out <= 64'd821107918729627811;
    11'd607: brom_out <= 64'd2749009972353655762;
    11'd608: brom_out <= 64'd3547627594494878621;
    11'd609: brom_out <= 64'd3136767173588347434;
    11'd610: brom_out <= 64'd1549287551893278911;
    11'd611: brom_out <= 64'd6579678929095156593;
    11'd612: brom_out <= 64'd57560180524151836;
    11'd613: brom_out <= 64'd8431525056773163324;
    11'd614: brom_out <= 64'd7831437647304356508;
    11'd615: brom_out <= 64'd25054386228368260;
    11'd616: brom_out <= 64'd5944864576936445287;
    11'd617: brom_out <= 64'd978720527126678484;
    11'd618: brom_out <= 64'd5078991997579173257;
    11'd619: brom_out <= 64'd5515184158531911546;
    11'd620: brom_out <= 64'd684639643803771175;
    11'd621: brom_out <= 64'd3281923340519708537;
    11'd622: brom_out <= 64'd3340259218302706899;
    11'd623: brom_out <= 64'd3591529433803820433;
    11'd624: brom_out <= 64'd2468663283803736374;
    11'd625: brom_out <= 64'd4585935009530136169;
    11'd626: brom_out <= 64'd5798824876843371582;
    11'd627: brom_out <= 64'd2212864360945965123;
    11'd628: brom_out <= 64'd1837680713908133646;
    11'd629: brom_out <= 64'd672919549451933827;
    11'd630: brom_out <= 64'd2036591841189774695;
    11'd631: brom_out <= 64'd6072046178105556475;
    11'd632: brom_out <= 64'd1178188298187125443;
    11'd633: brom_out <= 64'd5545686084666219710;
    11'd634: brom_out <= 64'd3110559949174149380;
    11'd635: brom_out <= 64'd1330381704714286085;
    11'd636: brom_out <= 64'd5873106135293020355;
    11'd637: brom_out <= 64'd1435120993511282705;
    11'd638: brom_out <= 64'd8803778985884906727;
    11'd639: brom_out <= 64'd6585546512385483974;
    11'd640: brom_out <= 64'd2991444385089030097;
    11'd641: brom_out <= 64'd6427097281726706628;
    11'd642: brom_out <= 64'd4183299227927339195;
    11'd643: brom_out <= 64'd3119079411128405209;
    11'd644: brom_out <= 64'd1122397655549924356;
    11'd645: brom_out <= 64'd5564951036314476973;
    11'd646: brom_out <= 64'd2527297775950676908;
    11'd647: brom_out <= 64'd3036875632463858834;
    11'd648: brom_out <= 64'd6281663284576107517;
    11'd649: brom_out <= 64'd4794722994419500598;
    11'd650: brom_out <= 64'd7533491753178725717;
    11'd651: brom_out <= 64'd8580562440646539131;
    11'd652: brom_out <= 64'd8697599446790123293;
    11'd653: brom_out <= 64'd5318448438505440257;
    11'd654: brom_out <= 64'd235142833563334451;
    11'd655: brom_out <= 64'd1078913570171309648;
    11'd656: brom_out <= 64'd8124953238658307565;
    11'd657: brom_out <= 64'd6514515671117556603;
    11'd658: brom_out <= 64'd5808776274764837854;
    11'd659: brom_out <= 64'd1737665055851572803;
    11'd660: brom_out <= 64'd4625294087119433729;
    11'd661: brom_out <= 64'd3148801124557623449;
    11'd662: brom_out <= 64'd75966845172534173;
    11'd663: brom_out <= 64'd1113248537812598346;
    11'd664: brom_out <= 64'd5782598045554155253;
    11'd665: brom_out <= 64'd1141036854004408858;
    11'd666: brom_out <= 64'd7870108581299121483;
    11'd667: brom_out <= 64'd4196968460687196785;
    11'd668: brom_out <= 64'd5991059833680697521;
    11'd669: brom_out <= 64'd4613903798598080436;
    11'd670: brom_out <= 64'd8100294372597586432;
    11'd671: brom_out <= 64'd3504473931275065124;
    11'd672: brom_out <= 64'd9166670786663116443;
    11'd673: brom_out <= 64'd5395617652967469222;
    11'd674: brom_out <= 64'd7083423175763586691;
    11'd675: brom_out <= 64'd7441158198174016671;
    11'd676: brom_out <= 64'd7173654840489607776;
    11'd677: brom_out <= 64'd8838718518559474163;
    11'd678: brom_out <= 64'd1947243181919420491;
    11'd679: brom_out <= 64'd3854484312171404456;
    11'd680: brom_out <= 64'd3115848091286679823;
    11'd681: brom_out <= 64'd8317588540207922448;
    11'd682: brom_out <= 64'd5226535173943436928;
    11'd683: brom_out <= 64'd3682273990606439039;
    11'd684: brom_out <= 64'd750361034814781007;
    11'd685: brom_out <= 64'd4397702267799328608;
    11'd686: brom_out <= 64'd3592198641247208794;
    11'd687: brom_out <= 64'd3433509905416311683;
    11'd688: brom_out <= 64'd5654726277541044038;
    11'd689: brom_out <= 64'd5083175541303528685;
    11'd690: brom_out <= 64'd4510264232516592952;
    11'd691: brom_out <= 64'd2931018764400806070;
    11'd692: brom_out <= 64'd5208814341045079371;
    11'd693: brom_out <= 64'd8312556079981528030;
    11'd694: brom_out <= 64'd5551115908770807940;
    11'd695: brom_out <= 64'd585096259269936048;
    11'd696: brom_out <= 64'd3558399091024426444;
    11'd697: brom_out <= 64'd4322711149969805068;
    11'd698: brom_out <= 64'd1491544262489362891;
    11'd699: brom_out <= 64'd6079977503648451335;
    11'd700: brom_out <= 64'd4764036910647300995;
    11'd701: brom_out <= 64'd1985994961055839280;
    11'd702: brom_out <= 64'd9197868711120196895;
    11'd703: brom_out <= 64'd6769971139694742693;
    11'd704: brom_out <= 64'd7646914504675205489;
    11'd705: brom_out <= 64'd8256294627998732981;
    11'd706: brom_out <= 64'd5713577346046003020;
    11'd707: brom_out <= 64'd1478979661686592040;
    11'd708: brom_out <= 64'd3065938557921374089;
    11'd709: brom_out <= 64'd2610367100111832212;
    11'd710: brom_out <= 64'd2744296939060575530;
    11'd711: brom_out <= 64'd3368411057424669635;
    11'd712: brom_out <= 64'd1555308162728177297;
    11'd713: brom_out <= 64'd4054013996166535507;
    11'd714: brom_out <= 64'd220088159844794260;
    11'd715: brom_out <= 64'd7976876523254192230;
    11'd716: brom_out <= 64'd6550225160897858344;
    11'd717: brom_out <= 64'd7892653319965062638;
    11'd718: brom_out <= 64'd5490294517849368108;
    11'd719: brom_out <= 64'd6199672516180526071;
    11'd720: brom_out <= 64'd2141707773911427712;
    11'd721: brom_out <= 64'd635855831193566106;
    11'd722: brom_out <= 64'd7593220218804307867;
    11'd723: brom_out <= 64'd8341925111666110475;
    11'd724: brom_out <= 64'd5418439566171715291;
    11'd725: brom_out <= 64'd8673620925411977753;
    11'd726: brom_out <= 64'd4249431574386262900;
    11'd727: brom_out <= 64'd2847404267546166357;
    11'd728: brom_out <= 64'd7010796944267998638;
    11'd729: brom_out <= 64'd3468411571066471426;
    11'd730: brom_out <= 64'd7135696680823117604;
    11'd731: brom_out <= 64'd6230035500739914156;
    11'd732: brom_out <= 64'd8692551628537520016;
    11'd733: brom_out <= 64'd8513076200388136183;
    11'd734: brom_out <= 64'd4824069180043442917;
    11'd735: brom_out <= 64'd1141842582310077908;
    11'd736: brom_out <= 64'd4393262027419573708;
    11'd737: brom_out <= 64'd3058650903359729066;
    11'd738: brom_out <= 64'd8893614490103508778;
    11'd739: brom_out <= 64'd7462328687096900295;
    11'd740: brom_out <= 64'd4159689793066360690;
    11'd741: brom_out <= 64'd6283534932199547339;
    11'd742: brom_out <= 64'd654752926994167022;
    11'd743: brom_out <= 64'd6628447066861725489;
    11'd744: brom_out <= 64'd4919595983980879989;
    11'd745: brom_out <= 64'd6301640391988730655;
    11'd746: brom_out <= 64'd2816403948006974041;
    11'd747: brom_out <= 64'd8969075915070151768;
    11'd748: brom_out <= 64'd4919750730687193807;
    11'd749: brom_out <= 64'd8694371873892844208;
    11'd750: brom_out <= 64'd4413826527383477878;
    11'd751: brom_out <= 64'd7030554445186196665;
    11'd752: brom_out <= 64'd5729951333194461427;
    11'd753: brom_out <= 64'd7978110531043641769;
    11'd754: brom_out <= 64'd8743332571195579934;
    11'd755: brom_out <= 64'd9129774312610320619;
    11'd756: brom_out <= 64'd2240289491309476277;
    11'd757: brom_out <= 64'd8440836487301065001;
    11'd758: brom_out <= 64'd2173356542276770935;
    11'd759: brom_out <= 64'd1755068967933061315;
    11'd760: brom_out <= 64'd1376701315345052441;
    11'd761: brom_out <= 64'd6593921752856366535;
    11'd762: brom_out <= 64'd3167756150689666531;
    11'd763: brom_out <= 64'd3784018163499518601;
    11'd764: brom_out <= 64'd5939667306004532036;
    11'd765: brom_out <= 64'd7427050020511569441;
    11'd766: brom_out <= 64'd2935114005611711057;
    11'd767: brom_out <= 64'd7692930341342185952;
    11'd768: brom_out <= 64'd3392617565049336557;
    11'd769: brom_out <= 64'd7131970059357333029;
    11'd770: brom_out <= 64'd2230049327513614869;
    11'd771: brom_out <= 64'd3854526127297200834;
    11'd772: brom_out <= 64'd7479147464852913991;
    11'd773: brom_out <= 64'd5742128143480654282;
    11'd774: brom_out <= 64'd7538107808473199530;
    11'd775: brom_out <= 64'd822715829145346347;
    11'd776: brom_out <= 64'd2263269548655216762;
    11'd777: brom_out <= 64'd3329822700088162495;
    11'd778: brom_out <= 64'd6798664954031634633;
    11'd779: brom_out <= 64'd4175560118002252921;
    11'd780: brom_out <= 64'd6982695801609760735;
    11'd781: brom_out <= 64'd6913663135607926584;
    11'd782: brom_out <= 64'd6068442745462420874;
    11'd783: brom_out <= 64'd2228552985412019277;
    11'd784: brom_out <= 64'd8216761589456164;
    11'd785: brom_out <= 64'd5266018003312504579;
    11'd786: brom_out <= 64'd9102413699342598757;
    11'd787: brom_out <= 64'd3580819943894297764;
    11'd788: brom_out <= 64'd6925371594294004533;
    11'd789: brom_out <= 64'd4784055077466289542;
    11'd790: brom_out <= 64'd1568136098664689522;
    11'd791: brom_out <= 64'd4419790281338715805;
    11'd792: brom_out <= 64'd8186964208105355814;
    11'd793: brom_out <= 64'd8817464271798224027;
    11'd794: brom_out <= 64'd1676869911627098617;
    11'd795: brom_out <= 64'd4401819749409430491;
    11'd796: brom_out <= 64'd6849437044168275747;
    11'd797: brom_out <= 64'd7286314464983170863;
    11'd798: brom_out <= 64'd8444867741212273661;
    11'd799: brom_out <= 64'd9151515973652221402;
    11'd800: brom_out <= 64'd5039744181953194803;
    11'd801: brom_out <= 64'd637799399688374479;
    11'd802: brom_out <= 64'd3468732936118861906;
    11'd803: brom_out <= 64'd2777986735042830839;
    11'd804: brom_out <= 64'd3064309850488305304;
    11'd805: brom_out <= 64'd4131185556170130308;
    11'd806: brom_out <= 64'd391518006782257654;
    11'd807: brom_out <= 64'd2051836413390839457;
    11'd808: brom_out <= 64'd5471972468712594632;
    11'd809: brom_out <= 64'd8595678383967341286;
    11'd810: brom_out <= 64'd8395167631823199941;
    11'd811: brom_out <= 64'd8907923421314590115;
    11'd812: brom_out <= 64'd6626178562688381462;
    11'd813: brom_out <= 64'd5769552562384596599;
    11'd814: brom_out <= 64'd9209536114756024834;
    11'd815: brom_out <= 64'd8947667063148711049;
    11'd816: brom_out <= 64'd1628906345678539120;
    11'd817: brom_out <= 64'd1544674224130596118;
    11'd818: brom_out <= 64'd4368700210148671551;
    11'd819: brom_out <= 64'd6319435406754674390;
    11'd820: brom_out <= 64'd7705829573832500897;
    11'd821: brom_out <= 64'd4677673593772524828;
    11'd822: brom_out <= 64'd4934228471949137670;
    11'd823: brom_out <= 64'd5511461520034253554;
    11'd824: brom_out <= 64'd3528090222809025860;
    11'd825: brom_out <= 64'd1607600945152906512;
    11'd826: brom_out <= 64'd1258669831230654444;
    11'd827: brom_out <= 64'd2170069437537526133;
    11'd828: brom_out <= 64'd8798316185508471405;
    11'd829: brom_out <= 64'd7183585907134239486;
    11'd830: brom_out <= 64'd6154077313509807261;
    11'd831: brom_out <= 64'd4955822627172985255;
    11'd832: brom_out <= 64'd1002059954001900696;
    11'd833: brom_out <= 64'd4687421323741025393;
    11'd834: brom_out <= 64'd2757773614559033666;
    11'd835: brom_out <= 64'd4725094368207763061;
    11'd836: brom_out <= 64'd1490887556607246244;
    11'd837: brom_out <= 64'd91987351604627050;
    11'd838: brom_out <= 64'd7104811893195087792;
    11'd839: brom_out <= 64'd7767226473893413332;
    11'd840: brom_out <= 64'd307156682351195017;
    11'd841: brom_out <= 64'd4898893176619253892;
    11'd842: brom_out <= 64'd8730278730941939396;
    11'd843: brom_out <= 64'd3005741243809146285;
    11'd844: brom_out <= 64'd3107918471259441615;
    11'd845: brom_out <= 64'd725251043603134492;
    11'd846: brom_out <= 64'd6460685242337216620;
    11'd847: brom_out <= 64'd5450767261026876886;
    11'd848: brom_out <= 64'd4836003352449041316;
    11'd849: brom_out <= 64'd956565536080223686;
    11'd850: brom_out <= 64'd8051296741047110195;
    11'd851: brom_out <= 64'd4077815017758764724;
    11'd852: brom_out <= 64'd2923414615723271043;
    11'd853: brom_out <= 64'd820027634638271577;
    11'd854: brom_out <= 64'd8026629062288902533;
    11'd855: brom_out <= 64'd2595667101902401433;
    11'd856: brom_out <= 64'd6436331060924184539;
    11'd857: brom_out <= 64'd5549270204663924183;
    11'd858: brom_out <= 64'd6733707155866364304;
    11'd859: brom_out <= 64'd546478178973529773;
    11'd860: brom_out <= 64'd1641922973023157952;
    11'd861: brom_out <= 64'd2003304190459111066;
    11'd862: brom_out <= 64'd4681773058202772675;
    11'd863: brom_out <= 64'd3404093846247594996;
    11'd864: brom_out <= 64'd9185509849420767578;
    11'd865: brom_out <= 64'd6282214430396223665;
    11'd866: brom_out <= 64'd6230952056441481807;
    11'd867: brom_out <= 64'd5651215856363377316;
    11'd868: brom_out <= 64'd1546731779372361302;
    11'd869: brom_out <= 64'd3758573853795653427;
    11'd870: brom_out <= 64'd1790792280522562723;
    11'd871: brom_out <= 64'd6760985867545539242;
    11'd872: brom_out <= 64'd7995675456769788758;
    11'd873: brom_out <= 64'd3111218648416961668;
    11'd874: brom_out <= 64'd198235807530720187;
    11'd875: brom_out <= 64'd5168690797098687629;
    11'd876: brom_out <= 64'd4849682055056439114;
    11'd877: brom_out <= 64'd1337980060505609637;
    11'd878: brom_out <= 64'd9160052455972965925;
    11'd879: brom_out <= 64'd6411251051681906994;
    11'd880: brom_out <= 64'd9003279055065478956;
    11'd881: brom_out <= 64'd3820044292411662612;
    11'd882: brom_out <= 64'd5011986474190685475;
    11'd883: brom_out <= 64'd8698260697543325537;
    11'd884: brom_out <= 64'd869826359180825983;
    11'd885: brom_out <= 64'd3445970765661623385;
    11'd886: brom_out <= 64'd6630229277550940928;
    11'd887: brom_out <= 64'd1664928300054969876;
    11'd888: brom_out <= 64'd1827606411485443129;
    11'd889: brom_out <= 64'd6181880917497703341;
    11'd890: brom_out <= 64'd6949147395764538964;
    11'd891: brom_out <= 64'd7253780654183843384;
    11'd892: brom_out <= 64'd7672998258368931866;
    11'd893: brom_out <= 64'd1950822828069733729;
    11'd894: brom_out <= 64'd7530731249570041776;
    11'd895: brom_out <= 64'd8631772682564570593;
    11'd896: brom_out <= 64'd699101306064864663;
    11'd897: brom_out <= 64'd7889711590670918676;
    11'd898: brom_out <= 64'd655123889431899961;
    11'd899: brom_out <= 64'd2126660867906687864;
    11'd900: brom_out <= 64'd8219959792660589692;
    11'd901: brom_out <= 64'd8551637415506572346;
    11'd902: brom_out <= 64'd8543830174923091154;
    11'd903: brom_out <= 64'd1435047781493708974;
    11'd904: brom_out <= 64'd5893272571222366297;
    11'd905: brom_out <= 64'd7027244046667068898;
    11'd906: brom_out <= 64'd2015889517693822068;
    11'd907: brom_out <= 64'd4971028798941293784;
    11'd908: brom_out <= 64'd4439925312673350003;
    11'd909: brom_out <= 64'd2408543357995828304;
    11'd910: brom_out <= 64'd4798734633597747276;
    11'd911: brom_out <= 64'd6781627562122407399;
    11'd912: brom_out <= 64'd69843017785227084;
    11'd913: brom_out <= 64'd4891530948138436991;
    11'd914: brom_out <= 64'd8247980103556855667;
    11'd915: brom_out <= 64'd2840283348677403338;
    11'd916: brom_out <= 64'd8225172405297280263;
    11'd917: brom_out <= 64'd7450817543983322844;
    11'd918: brom_out <= 64'd976868090527140556;
    11'd919: brom_out <= 64'd6363705655307338806;
    11'd920: brom_out <= 64'd7645071031480098655;
    11'd921: brom_out <= 64'd3868531777045828691;
    11'd922: brom_out <= 64'd5140288024937627165;
    11'd923: brom_out <= 64'd4538780524597464161;
    11'd924: brom_out <= 64'd5173422508798334624;
    11'd925: brom_out <= 64'd5708860785940369427;
    11'd926: brom_out <= 64'd2600298912569494844;
    11'd927: brom_out <= 64'd6716916671807146392;
    11'd928: brom_out <= 64'd7923677684682802987;
    11'd929: brom_out <= 64'd3815011943812575350;
    11'd930: brom_out <= 64'd2275953281661646751;
    11'd931: brom_out <= 64'd5745260692505968145;
    11'd932: brom_out <= 64'd2139689406997953411;
    11'd933: brom_out <= 64'd8748419681862114146;
    11'd934: brom_out <= 64'd3729764982569583119;
    11'd935: brom_out <= 64'd1674345919730951813;
    11'd936: brom_out <= 64'd375356035198548383;
    11'd937: brom_out <= 64'd1373369117410510866;
    11'd938: brom_out <= 64'd4961919869715327681;
    11'd939: brom_out <= 64'd9052054262515000354;
    11'd940: brom_out <= 64'd511527761999251354;
    11'd941: brom_out <= 64'd3482983880212475854;
    11'd942: brom_out <= 64'd5412893724914022449;
    11'd943: brom_out <= 64'd5032214272686406166;
    11'd944: brom_out <= 64'd5126845061066175356;
    11'd945: brom_out <= 64'd7984550382453767596;
    11'd946: brom_out <= 64'd6181066534637459237;
    11'd947: brom_out <= 64'd8680510475920407927;
    11'd948: brom_out <= 64'd9162350688835803463;
    11'd949: brom_out <= 64'd1414658525045134853;
    11'd950: brom_out <= 64'd841949363898762459;
    11'd951: brom_out <= 64'd486400348447004409;
    11'd952: brom_out <= 64'd796180145389681740;
    11'd953: brom_out <= 64'd8371723383654335520;
    11'd954: brom_out <= 64'd6881112568257936145;
    11'd955: brom_out <= 64'd8219861536954301229;
    11'd956: brom_out <= 64'd4119508171639317112;
    11'd957: brom_out <= 64'd2072885801364544572;
    11'd958: brom_out <= 64'd4523573697502160143;
    11'd959: brom_out <= 64'd9096591304164137574;
    11'd960: brom_out <= 64'd1670791095363685175;
    11'd961: brom_out <= 64'd3613147540994151386;
    11'd962: brom_out <= 64'd6268445540391799960;
    11'd963: brom_out <= 64'd333801395018402419;
    11'd964: brom_out <= 64'd5989914729659460893;
    11'd965: brom_out <= 64'd5421197279853390596;
    11'd966: brom_out <= 64'd8498706274306490892;
    11'd967: brom_out <= 64'd7292703967224865486;
    11'd968: brom_out <= 64'd3280526131456603436;
    11'd969: brom_out <= 64'd291195603844344417;
    11'd970: brom_out <= 64'd881381962624186811;
    11'd971: brom_out <= 64'd2351202851047628420;
    11'd972: brom_out <= 64'd3615127351505505023;
    11'd973: brom_out <= 64'd6062993788722341892;
    11'd974: brom_out <= 64'd6148609810148795929;
    11'd975: brom_out <= 64'd599730283692523374;
    11'd976: brom_out <= 64'd8823464365455855293;
    11'd977: brom_out <= 64'd5749262411298578370;
    11'd978: brom_out <= 64'd5139097896322553033;
    11'd979: brom_out <= 64'd8165494333656525134;
    11'd980: brom_out <= 64'd5003529372930301250;
    11'd981: brom_out <= 64'd6319980041019054251;
    11'd982: brom_out <= 64'd3363566323249637328;
    11'd983: brom_out <= 64'd5252122029312962963;
    11'd984: brom_out <= 64'd8323983203612776937;
    11'd985: brom_out <= 64'd2040235830658135393;
    11'd986: brom_out <= 64'd3740576396473059045;
    11'd987: brom_out <= 64'd3289458284692175700;
    11'd988: brom_out <= 64'd5423351720389833865;
    11'd989: brom_out <= 64'd2497038050456785463;
    11'd990: brom_out <= 64'd5408302969401217960;
    11'd991: brom_out <= 64'd7848005646647114461;
    11'd992: brom_out <= 64'd228503451388919711;
    11'd993: brom_out <= 64'd2939264214977633037;
    11'd994: brom_out <= 64'd6913883903315781469;
    11'd995: brom_out <= 64'd3506647722126204218;
    11'd996: brom_out <= 64'd498968785704607628;
    11'd997: brom_out <= 64'd911760100456784026;
    11'd998: brom_out <= 64'd3083280881619226755;
    11'd999: brom_out <= 64'd4628098658155976042;
    11'd1000: brom_out <= 64'd7002130558985726630;
    11'd1001: brom_out <= 64'd2804463966393397031;
    11'd1002: brom_out <= 64'd3016980039216328962;
    11'd1003: brom_out <= 64'd7857926944957203380;
    11'd1004: brom_out <= 64'd7471415495952780188;
    11'd1005: brom_out <= 64'd713405409942497823;
    11'd1006: brom_out <= 64'd9117660520541870682;
    11'd1007: brom_out <= 64'd333363560357025169;
    11'd1008: brom_out <= 64'd700730835196570872;
    11'd1009: brom_out <= 64'd646297118098278772;
    11'd1010: brom_out <= 64'd7087203385146507098;
    11'd1011: brom_out <= 64'd2133757072145401712;
    11'd1012: brom_out <= 64'd8584995141337045279;
    11'd1013: brom_out <= 64'd830325714398867404;
    11'd1014: brom_out <= 64'd6918964554399920495;
    11'd1015: brom_out <= 64'd8758553949588800273;
    11'd1016: brom_out <= 64'd2113561489472542490;
    11'd1017: brom_out <= 64'd4130478540001382116;
    11'd1018: brom_out <= 64'd3835383961103183096;
    11'd1019: brom_out <= 64'd2997007021939187347;
    11'd1020: brom_out <= 64'd7269045898348823146;
    11'd1021: brom_out <= 64'd3031303078308718036;
    11'd1022: brom_out <= 64'd8634110784643349010;
    11'd1023: brom_out <= 64'd4803548634770013292;
    default: brom_out <= 64'h1;
    endcase
end

generate
    if(DELAY == 1) begin
        assign b = brom_out;
    end
endgenerate

endmodule

//-------------------------------------------------------------------------------------------------

module tw_rom_11
#(
    parameter LOGN  = 11,
    parameter LOGQ  = 64,
    parameter DELAY = 1,
    parameter STAGE = 1
)(
    input            clk,
    input [LOGN-1:0] raddr,
    output[LOGQ-1:0] b
);

(* ram_style = "block" *)
reg [LOGQ-1:0] brom_out, brom_out2;

always @(posedge clk) begin
    case(raddr[STAGE-1:0])
    12'd0: brom_out <= 64'd9223372036854251519;
    12'd1: brom_out <= 64'd1102913100553729005;
    12'd2: brom_out <= 64'd6012871302989280084;
    12'd3: brom_out <= 64'd1527009950824020455;
    12'd4: brom_out <= 64'd7605493872853681221;
    12'd5: brom_out <= 64'd331705278823141530;
    12'd6: brom_out <= 64'd3127052517479868225;
    12'd7: brom_out <= 64'd4972921688478999892;
    12'd8: brom_out <= 64'd1299456045732977605;
    12'd9: brom_out <= 64'd5667686056105230206;
    12'd10: brom_out <= 64'd9150256334426485369;
    12'd11: brom_out <= 64'd7706649108346001651;
    12'd12: brom_out <= 64'd8213948439719346069;
    12'd13: brom_out <= 64'd7172243811045393643;
    12'd14: brom_out <= 64'd6825597430088558793;
    12'd15: brom_out <= 64'd3948706956136277229;
    12'd16: brom_out <= 64'd269998454485676360;
    12'd17: brom_out <= 64'd7325184581455921607;
    12'd18: brom_out <= 64'd2564423744727517704;
    12'd19: brom_out <= 64'd6682290189906599342;
    12'd20: brom_out <= 64'd7934371085285641861;
    12'd21: brom_out <= 64'd3326814094761790440;
    12'd22: brom_out <= 64'd7153207102067290344;
    12'd23: brom_out <= 64'd5020486994570292715;
    12'd24: brom_out <= 64'd9033387621081412018;
    12'd25: brom_out <= 64'd6205137676891788173;
    12'd26: brom_out <= 64'd3293074636399430213;
    12'd27: brom_out <= 64'd1238696719636161094;
    12'd28: brom_out <= 64'd4765886196678305331;
    12'd29: brom_out <= 64'd6624943704144324919;
    12'd30: brom_out <= 64'd5112583091541522973;
    12'd31: brom_out <= 64'd4373906864111961192;
    12'd32: brom_out <= 64'd6984365454624050605;
    12'd33: brom_out <= 64'd344548888781770986;
    12'd34: brom_out <= 64'd2273617654662494576;
    12'd35: brom_out <= 64'd1572845108645829558;
    12'd36: brom_out <= 64'd2123066514724381883;
    12'd37: brom_out <= 64'd8549720275696150946;
    12'd38: brom_out <= 64'd2567313654253520317;
    12'd39: brom_out <= 64'd9089944754788158967;
    12'd40: brom_out <= 64'd810060818546034655;
    12'd41: brom_out <= 64'd3777600355184077437;
    12'd42: brom_out <= 64'd6588969549873072984;
    12'd43: brom_out <= 64'd5984646794750834878;
    12'd44: brom_out <= 64'd8581206737579399620;
    12'd45: brom_out <= 64'd331112463124969936;
    12'd46: brom_out <= 64'd7820318430984191122;
    12'd47: brom_out <= 64'd8404649338598950687;
    12'd48: brom_out <= 64'd5653377166457707394;
    12'd49: brom_out <= 64'd3839782310825792117;
    12'd50: brom_out <= 64'd2934009396408142147;
    12'd51: brom_out <= 64'd6615922998039242763;
    12'd52: brom_out <= 64'd2299841007653134372;
    12'd53: brom_out <= 64'd5069310872664059544;
    12'd54: brom_out <= 64'd1287674294028378649;
    12'd55: brom_out <= 64'd543826894803705978;
    12'd56: brom_out <= 64'd8914698016797979130;
    12'd57: brom_out <= 64'd3169786119895682072;
    12'd58: brom_out <= 64'd4290018412507268451;
    12'd59: brom_out <= 64'd957479872005410401;
    12'd60: brom_out <= 64'd5779395201958353378;
    12'd61: brom_out <= 64'd7758685808708086097;
    12'd62: brom_out <= 64'd8710174058585331351;
    12'd63: brom_out <= 64'd5596293620407173703;
    12'd64: brom_out <= 64'd8706294438413809553;
    12'd65: brom_out <= 64'd3702518847184112432;
    12'd66: brom_out <= 64'd6756792246403704650;
    12'd67: brom_out <= 64'd5445518581501875667;
    12'd68: brom_out <= 64'd2509796222201502174;
    12'd69: brom_out <= 64'd494274216377378736;
    12'd70: brom_out <= 64'd1467033842096743702;
    12'd71: brom_out <= 64'd1476514077331314976;
    12'd72: brom_out <= 64'd1984480336129885140;
    12'd73: brom_out <= 64'd819099372979029972;
    12'd74: brom_out <= 64'd5411415188401616703;
    12'd75: brom_out <= 64'd1757503418561083295;
    12'd76: brom_out <= 64'd7152306933764292478;
    12'd77: brom_out <= 64'd5208933208073689448;
    12'd78: brom_out <= 64'd8367416970837404480;
    12'd79: brom_out <= 64'd5002790962071147126;
    12'd80: brom_out <= 64'd6626061600160634657;
    12'd81: brom_out <= 64'd7849000344767537809;
    12'd82: brom_out <= 64'd1408687539684857079;
    12'd83: brom_out <= 64'd3614648718488622517;
    12'd84: brom_out <= 64'd4332795524147639451;
    12'd85: brom_out <= 64'd4416538491726633807;
    12'd86: brom_out <= 64'd6891504871357446422;
    12'd87: brom_out <= 64'd4987120826118502355;
    12'd88: brom_out <= 64'd6375267241083926885;
    12'd89: brom_out <= 64'd5281767851388166670;
    12'd90: brom_out <= 64'd7586867602903602858;
    12'd91: brom_out <= 64'd4765428132147807493;
    12'd92: brom_out <= 64'd792297214988562254;
    12'd93: brom_out <= 64'd5290510743141442020;
    12'd94: brom_out <= 64'd7058677087284092182;
    12'd95: brom_out <= 64'd1674291621165505607;
    12'd96: brom_out <= 64'd6158485483849164736;
    12'd97: brom_out <= 64'd5160493589408218780;
    12'd98: brom_out <= 64'd5266916899250488660;
    12'd99: brom_out <= 64'd2125871470203471318;
    12'd100: brom_out <= 64'd1966154900029444318;
    12'd101: brom_out <= 64'd7970308623799195545;
    12'd102: brom_out <= 64'd1215003878949612048;
    12'd103: brom_out <= 64'd6376806131588433218;
    12'd104: brom_out <= 64'd2808688244394002011;
    12'd105: brom_out <= 64'd1857577982111137819;
    12'd106: brom_out <= 64'd3851039626226392450;
    12'd107: brom_out <= 64'd6186730927293561609;
    12'd108: brom_out <= 64'd7902540812321798218;
    12'd109: brom_out <= 64'd7685174008941584275;
    12'd110: brom_out <= 64'd6004430279489338680;
    12'd111: brom_out <= 64'd5215512869855517538;
    12'd112: brom_out <= 64'd7345482494331839697;
    12'd113: brom_out <= 64'd453811032764871892;
    12'd114: brom_out <= 64'd4218632253198916038;
    12'd115: brom_out <= 64'd4326695183155906556;
    12'd116: brom_out <= 64'd299894953115934099;
    12'd117: brom_out <= 64'd8426041380979419904;
    12'd118: brom_out <= 64'd1821424608084578998;
    12'd119: brom_out <= 64'd4350436591725259429;
    12'd120: brom_out <= 64'd8037037384829722617;
    12'd121: brom_out <= 64'd222767951529780175;
    12'd122: brom_out <= 64'd4110036900460384796;
    12'd123: brom_out <= 64'd8106152487619506999;
    12'd124: brom_out <= 64'd9104612624170912214;
    12'd125: brom_out <= 64'd4481386419402181357;
    12'd126: brom_out <= 64'd1547693224024900634;
    12'd127: brom_out <= 64'd8674474176990565409;
    12'd128: brom_out <= 64'd5917339183240377480;
    12'd129: brom_out <= 64'd2038520525822259048;
    12'd130: brom_out <= 64'd8498480881154740865;
    12'd131: brom_out <= 64'd5587791659679814202;
    12'd132: brom_out <= 64'd4392041727794040139;
    12'd133: brom_out <= 64'd4507188278956917814;
    12'd134: brom_out <= 64'd6475240946856553091;
    12'd135: brom_out <= 64'd2922269551779043038;
    12'd136: brom_out <= 64'd3561119328844693546;
    12'd137: brom_out <= 64'd1625945569422476240;
    12'd138: brom_out <= 64'd5569609541362591627;
    12'd139: brom_out <= 64'd5345829616181158893;
    12'd140: brom_out <= 64'd2908884142996516879;
    12'd141: brom_out <= 64'd5267269215936573461;
    12'd142: brom_out <= 64'd3495906847793555496;
    12'd143: brom_out <= 64'd8152988480412639353;
    12'd144: brom_out <= 64'd8174323033676948403;
    12'd145: brom_out <= 64'd418688512246794328;
    12'd146: brom_out <= 64'd8346874721972884401;
    12'd147: brom_out <= 64'd8897437151834909042;
    12'd148: brom_out <= 64'd7153542761736184733;
    12'd149: brom_out <= 64'd4599926363795950470;
    12'd150: brom_out <= 64'd9036614214691043214;
    12'd151: brom_out <= 64'd6430137174595182183;
    12'd152: brom_out <= 64'd2319035647868930894;
    12'd153: brom_out <= 64'd8927043086982599750;
    12'd154: brom_out <= 64'd1331680507007219705;
    12'd155: brom_out <= 64'd8668330478160946558;
    12'd156: brom_out <= 64'd5900439431409958858;
    12'd157: brom_out <= 64'd6037508690161556393;
    12'd158: brom_out <= 64'd8944063972887106670;
    12'd159: brom_out <= 64'd991733121096816246;
    12'd160: brom_out <= 64'd3950921523134993168;
    12'd161: brom_out <= 64'd5945019363494978713;
    12'd162: brom_out <= 64'd2884516234218684811;
    12'd163: brom_out <= 64'd4374432210238539416;
    12'd164: brom_out <= 64'd2162992210110465427;
    12'd165: brom_out <= 64'd5227741310768365469;
    12'd166: brom_out <= 64'd7920402332462387511;
    12'd167: brom_out <= 64'd2473325997743944052;
    12'd168: brom_out <= 64'd3531419639158455240;
    12'd169: brom_out <= 64'd328762820884200268;
    12'd170: brom_out <= 64'd7396774219033937672;
    12'd171: brom_out <= 64'd3958484914374424336;
    12'd172: brom_out <= 64'd6297866057014224030;
    12'd173: brom_out <= 64'd2887841837436318313;
    12'd174: brom_out <= 64'd1188483528343374386;
    12'd175: brom_out <= 64'd8745925251385352737;
    12'd176: brom_out <= 64'd4573453364429337213;
    12'd177: brom_out <= 64'd6432855811330329932;
    12'd178: brom_out <= 64'd6252329300465472480;
    12'd179: brom_out <= 64'd4625169900183292974;
    12'd180: brom_out <= 64'd1287149587930120656;
    12'd181: brom_out <= 64'd4975661477061904853;
    12'd182: brom_out <= 64'd5698207036020272794;
    12'd183: brom_out <= 64'd2851129277900631036;
    12'd184: brom_out <= 64'd3367056065757602806;
    12'd185: brom_out <= 64'd2387994583949301874;
    12'd186: brom_out <= 64'd118243567567768095;
    12'd187: brom_out <= 64'd3670854517306604647;
    12'd188: brom_out <= 64'd3883460632785907410;
    12'd189: brom_out <= 64'd9058002763678952859;
    12'd190: brom_out <= 64'd4486934250525894693;
    12'd191: brom_out <= 64'd7138994063059429231;
    12'd192: brom_out <= 64'd4110363107264655732;
    12'd193: brom_out <= 64'd1189672448575511328;
    12'd194: brom_out <= 64'd4514892859148397044;
    12'd195: brom_out <= 64'd4047332604529772758;
    12'd196: brom_out <= 64'd5549948750888088698;
    12'd197: brom_out <= 64'd2103746687090801379;
    12'd198: brom_out <= 64'd2943321537520600659;
    12'd199: brom_out <= 64'd13677257000361224;
    12'd200: brom_out <= 64'd5233426006749936404;
    12'd201: brom_out <= 64'd2916236583736325519;
    12'd202: brom_out <= 64'd5747717726212286166;
    12'd203: brom_out <= 64'd7181474872531538448;
    12'd204: brom_out <= 64'd7125634071680409905;
    12'd205: brom_out <= 64'd3520800072367565818;
    12'd206: brom_out <= 64'd4614122134803297477;
    12'd207: brom_out <= 64'd4254624995020049834;
    12'd208: brom_out <= 64'd8070303386396255336;
    12'd209: brom_out <= 64'd3900996048308082675;
    12'd210: brom_out <= 64'd8117367890929318445;
    12'd211: brom_out <= 64'd7126809288095688532;
    12'd212: brom_out <= 64'd4346701462512900589;
    12'd213: brom_out <= 64'd5226018621464696967;
    12'd214: brom_out <= 64'd7783606212229745263;
    12'd215: brom_out <= 64'd3590495931749359103;
    12'd216: brom_out <= 64'd5682374489572555945;
    12'd217: brom_out <= 64'd5025424451158582242;
    12'd218: brom_out <= 64'd880050980480071141;
    12'd219: brom_out <= 64'd3219436865258312315;
    12'd220: brom_out <= 64'd173114810237193158;
    12'd221: brom_out <= 64'd224320552559350026;
    12'd222: brom_out <= 64'd5314247580215590840;
    12'd223: brom_out <= 64'd7186500760229875053;
    12'd224: brom_out <= 64'd2194362728065833183;
    12'd225: brom_out <= 64'd7500931859087234329;
    12'd226: brom_out <= 64'd7403262497201993765;
    12'd227: brom_out <= 64'd3907478483338414094;
    12'd228: brom_out <= 64'd401958369407258982;
    12'd229: brom_out <= 64'd6887711032745255742;
    12'd230: brom_out <= 64'd4151717614504932492;
    12'd231: brom_out <= 64'd6460853876874714811;
    12'd232: brom_out <= 64'd240070673848085803;
    12'd233: brom_out <= 64'd7333325376921592110;
    12'd234: brom_out <= 64'd4057166001169818856;
    12'd235: brom_out <= 64'd2683430372073479744;
    12'd236: brom_out <= 64'd1427846036265206780;
    12'd237: brom_out <= 64'd765045619723753688;
    12'd238: brom_out <= 64'd5295131112655049137;
    12'd239: brom_out <= 64'd7386813248718022410;
    12'd240: brom_out <= 64'd6564530672913887453;
    12'd241: brom_out <= 64'd7103911473611199541;
    12'd242: brom_out <= 64'd3866632472152804465;
    12'd243: brom_out <= 64'd2104670626740145188;
    12'd244: brom_out <= 64'd3098083654159802861;
    12'd245: brom_out <= 64'd2203451223094322762;
    12'd246: brom_out <= 64'd3063481684957609078;
    12'd247: brom_out <= 64'd7972835908627627311;
    12'd248: brom_out <= 64'd1907082839763808740;
    12'd249: brom_out <= 64'd7686709619505464880;
    12'd250: brom_out <= 64'd1468430662791236228;
    12'd251: brom_out <= 64'd8995510598615158165;
    12'd252: brom_out <= 64'd3031844387819961827;
    12'd253: brom_out <= 64'd4390718853010686896;
    12'd254: brom_out <= 64'd1396316958451531348;
    12'd255: brom_out <= 64'd1680679157528580243;
    12'd256: brom_out <= 64'd2881966912403406253;
    12'd257: brom_out <= 64'd2801867022993033546;
    12'd258: brom_out <= 64'd9146187461299601623;
    12'd259: brom_out <= 64'd2918757492399093761;
    12'd260: brom_out <= 64'd2925409531261716840;
    12'd261: brom_out <= 64'd9125104620207024390;
    12'd262: brom_out <= 64'd4304180803912282259;
    12'd263: brom_out <= 64'd7003030798630255435;
    12'd264: brom_out <= 64'd8852621130615879035;
    12'd265: brom_out <= 64'd7303964566607951423;
    12'd266: brom_out <= 64'd4848840577486999766;
    12'd267: brom_out <= 64'd4368601964820485477;
    12'd268: brom_out <= 64'd270496797777326527;
    12'd269: brom_out <= 64'd5923984013916025162;
    12'd270: brom_out <= 64'd6083010805285052716;
    12'd271: brom_out <= 64'd1194702245926272972;
    12'd272: brom_out <= 64'd1219064800028085468;
    12'd273: brom_out <= 64'd1779228674047657867;
    12'd274: brom_out <= 64'd6306667576969932326;
    12'd275: brom_out <= 64'd6435347175821900655;
    12'd276: brom_out <= 64'd543577740076728061;
    12'd277: brom_out <= 64'd4863463436130572984;
    12'd278: brom_out <= 64'd4091222591604623441;
    12'd279: brom_out <= 64'd6904042720651947488;
    12'd280: brom_out <= 64'd1865389637899575391;
    12'd281: brom_out <= 64'd3873586375647389700;
    12'd282: brom_out <= 64'd2862891865227566885;
    12'd283: brom_out <= 64'd8216846839876223100;
    12'd284: brom_out <= 64'd7923340214113792441;
    12'd285: brom_out <= 64'd4899537041491779759;
    12'd286: brom_out <= 64'd4822434129781452362;
    12'd287: brom_out <= 64'd3405667996999341347;
    12'd288: brom_out <= 64'd735439083491420630;
    12'd289: brom_out <= 64'd4414035617291553258;
    12'd290: brom_out <= 64'd8701208384429075876;
    12'd291: brom_out <= 64'd1642318664855664016;
    12'd292: brom_out <= 64'd5356334136853441455;
    12'd293: brom_out <= 64'd339881140317908839;
    12'd294: brom_out <= 64'd2004505146951275140;
    12'd295: brom_out <= 64'd6254333483692308558;
    12'd296: brom_out <= 64'd4936662293846854616;
    12'd297: brom_out <= 64'd3773506948494418480;
    12'd298: brom_out <= 64'd695669619354178199;
    12'd299: brom_out <= 64'd7508137942481891379;
    12'd300: brom_out <= 64'd5689831925774807956;
    12'd301: brom_out <= 64'd7801453391915490838;
    12'd302: brom_out <= 64'd1189038338221773258;
    12'd303: brom_out <= 64'd2642030319808362412;
    12'd304: brom_out <= 64'd544940125055465581;
    12'd305: brom_out <= 64'd8988022062613589533;
    12'd306: brom_out <= 64'd2331992164875830888;
    12'd307: brom_out <= 64'd3496349151480100481;
    12'd308: brom_out <= 64'd1297536695137410486;
    12'd309: brom_out <= 64'd5215432719681743341;
    12'd310: brom_out <= 64'd4174433604295068968;
    12'd311: brom_out <= 64'd4108995439916808286;
    12'd312: brom_out <= 64'd1845447672304840611;
    12'd313: brom_out <= 64'd8580338531199479822;
    12'd314: brom_out <= 64'd7530083780768442237;
    12'd315: brom_out <= 64'd8594835602539730064;
    12'd316: brom_out <= 64'd2182902326656347159;
    12'd317: brom_out <= 64'd3010982391224114088;
    12'd318: brom_out <= 64'd7697402264257745017;
    12'd319: brom_out <= 64'd8308116381684268102;
    12'd320: brom_out <= 64'd1624553938728686361;
    12'd321: brom_out <= 64'd4369822744919577129;
    12'd322: brom_out <= 64'd2235543617824736075;
    12'd323: brom_out <= 64'd7392630178923620229;
    12'd324: brom_out <= 64'd3012117742719754636;
    12'd325: brom_out <= 64'd5773608516567397090;
    12'd326: brom_out <= 64'd8395034085139528506;
    12'd327: brom_out <= 64'd6184511926724241706;
    12'd328: brom_out <= 64'd3586995478868233709;
    12'd329: brom_out <= 64'd4100239665487453604;
    12'd330: brom_out <= 64'd5121098992128955161;
    12'd331: brom_out <= 64'd6197181412830849464;
    12'd332: brom_out <= 64'd2057313745147478637;
    12'd333: brom_out <= 64'd7157945453815143715;
    12'd334: brom_out <= 64'd5160625525529957528;
    12'd335: brom_out <= 64'd1656556474370501420;
    12'd336: brom_out <= 64'd2926075365041679386;
    12'd337: brom_out <= 64'd1331624447098205033;
    12'd338: brom_out <= 64'd3516066647433260551;
    12'd339: brom_out <= 64'd3460988223109260373;
    12'd340: brom_out <= 64'd7993764406966422987;
    12'd341: brom_out <= 64'd3517922268454075034;
    12'd342: brom_out <= 64'd8037258735659770483;
    12'd343: brom_out <= 64'd7433176994362088473;
    12'd344: brom_out <= 64'd5712154480457087476;
    12'd345: brom_out <= 64'd5844731795589899787;
    12'd346: brom_out <= 64'd3018928514936204385;
    12'd347: brom_out <= 64'd4925083064398185451;
    12'd348: brom_out <= 64'd3479065458090349436;
    12'd349: brom_out <= 64'd2073611639215184113;
    12'd350: brom_out <= 64'd1585371721068583241;
    12'd351: brom_out <= 64'd4523172126112293441;
    12'd352: brom_out <= 64'd5875474638474206446;
    12'd353: brom_out <= 64'd3827692355908478929;
    12'd354: brom_out <= 64'd4515128673629883118;
    12'd355: brom_out <= 64'd8381509481982198757;
    12'd356: brom_out <= 64'd6548403254923287631;
    12'd357: brom_out <= 64'd8471785160522617325;
    12'd358: brom_out <= 64'd4752592209480917425;
    12'd359: brom_out <= 64'd8890166281502929697;
    12'd360: brom_out <= 64'd7289325041362829578;
    12'd361: brom_out <= 64'd3147501462716504700;
    12'd362: brom_out <= 64'd6185725345812273456;
    12'd363: brom_out <= 64'd3785970388161490303;
    12'd364: brom_out <= 64'd1785088414017673288;
    12'd365: brom_out <= 64'd8308285389689614985;
    12'd366: brom_out <= 64'd4798463378767722612;
    12'd367: brom_out <= 64'd3145699679273069605;
    12'd368: brom_out <= 64'd6222003843073247882;
    12'd369: brom_out <= 64'd1352173756344525495;
    12'd370: brom_out <= 64'd3324417521285869935;
    12'd371: brom_out <= 64'd3261813778574482554;
    12'd372: brom_out <= 64'd1990992240235617717;
    12'd373: brom_out <= 64'd2475140240274188043;
    12'd374: brom_out <= 64'd8528027318223251457;
    12'd375: brom_out <= 64'd8728287108636576294;
    12'd376: brom_out <= 64'd616529505270125954;
    12'd377: brom_out <= 64'd6619360377626727946;
    12'd378: brom_out <= 64'd1960716502804548672;
    12'd379: brom_out <= 64'd1296572473256973960;
    12'd380: brom_out <= 64'd4535501105232824056;
    12'd381: brom_out <= 64'd4682354897801007425;
    12'd382: brom_out <= 64'd2293080637268173952;
    12'd383: brom_out <= 64'd1549853121982486025;
    12'd384: brom_out <= 64'd7147821265559899415;
    12'd385: brom_out <= 64'd7574768217639654355;
    12'd386: brom_out <= 64'd8249092968287330570;
    12'd387: brom_out <= 64'd4643101887081870411;
    12'd388: brom_out <= 64'd1598994064067110291;
    12'd389: brom_out <= 64'd3050172956909809872;
    12'd390: brom_out <= 64'd6446311831687328438;
    12'd391: brom_out <= 64'd39054179753570328;
    12'd392: brom_out <= 64'd3149227341269420724;
    12'd393: brom_out <= 64'd1687881817758787752;
    12'd394: brom_out <= 64'd2519301650103661960;
    12'd395: brom_out <= 64'd61829322818278264;
    12'd396: brom_out <= 64'd904660340594613265;
    12'd397: brom_out <= 64'd998185447878790241;
    12'd398: brom_out <= 64'd3412151563337741352;
    12'd399: brom_out <= 64'd1014540976961417578;
    12'd400: brom_out <= 64'd4717392765204693644;
    12'd401: brom_out <= 64'd7248112848643534511;
    12'd402: brom_out <= 64'd865268308687100412;
    12'd403: brom_out <= 64'd6806940559200776408;
    12'd404: brom_out <= 64'd4359339040815035935;
    12'd405: brom_out <= 64'd2683991028645697880;
    12'd406: brom_out <= 64'd5458238346969861276;
    12'd407: brom_out <= 64'd1552474800957627860;
    12'd408: brom_out <= 64'd4312120720500409507;
    12'd409: brom_out <= 64'd5105669458685259425;
    12'd410: brom_out <= 64'd3241756220799506222;
    12'd411: brom_out <= 64'd5888155221788109374;
    12'd412: brom_out <= 64'd749037117208255733;
    12'd413: brom_out <= 64'd7293739831641998651;
    12'd414: brom_out <= 64'd8021309328199436730;
    12'd415: brom_out <= 64'd964260620430079549;
    12'd416: brom_out <= 64'd8826561644056073004;
    12'd417: brom_out <= 64'd4215582806609882491;
    12'd418: brom_out <= 64'd6492936536869808625;
    12'd419: brom_out <= 64'd8013752277862596731;
    12'd420: brom_out <= 64'd6153283181782085767;
    12'd421: brom_out <= 64'd8527813612084473546;
    12'd422: brom_out <= 64'd3042490808619695370;
    12'd423: brom_out <= 64'd7318487377759942214;
    12'd424: brom_out <= 64'd7048641871031816;
    12'd425: brom_out <= 64'd2602683653691326026;
    12'd426: brom_out <= 64'd6938251047297990533;
    12'd427: brom_out <= 64'd6146878404415362577;
    12'd428: brom_out <= 64'd3017602207931310620;
    12'd429: brom_out <= 64'd8008558357275281990;
    12'd430: brom_out <= 64'd6526255316566008010;
    12'd431: brom_out <= 64'd3949377814362547728;
    12'd432: brom_out <= 64'd3526492789053904424;
    12'd433: brom_out <= 64'd5738954251284061668;
    12'd434: brom_out <= 64'd1097341705165972594;
    12'd435: brom_out <= 64'd4059622768511913746;
    12'd436: brom_out <= 64'd489108130890476637;
    12'd437: brom_out <= 64'd6623537519035813176;
    12'd438: brom_out <= 64'd9168100354083393324;
    12'd439: brom_out <= 64'd1585427658453945272;
    12'd440: brom_out <= 64'd5311697839062869272;
    12'd441: brom_out <= 64'd5868434889645250855;
    12'd442: brom_out <= 64'd3754010688254048597;
    12'd443: brom_out <= 64'd1345532271632170682;
    12'd444: brom_out <= 64'd7009454947613216741;
    12'd445: brom_out <= 64'd2426069432682723438;
    12'd446: brom_out <= 64'd1722163249877292090;
    12'd447: brom_out <= 64'd7442965855326153148;
    12'd448: brom_out <= 64'd3044098306375364542;
    12'd449: brom_out <= 64'd1203939852511973662;
    12'd450: brom_out <= 64'd3652792854953481228;
    12'd451: brom_out <= 64'd6605244667463568635;
    12'd452: brom_out <= 64'd967392942188980461;
    12'd453: brom_out <= 64'd8216179491009474193;
    12'd454: brom_out <= 64'd494499881005363032;
    12'd455: brom_out <= 64'd3238882406020454937;
    12'd456: brom_out <= 64'd7940586545958498989;
    12'd457: brom_out <= 64'd4875826095999072140;
    12'd458: brom_out <= 64'd5108575401283476645;
    12'd459: brom_out <= 64'd143958327396720651;
    12'd460: brom_out <= 64'd8888883322669091370;
    12'd461: brom_out <= 64'd1006312549628104935;
    12'd462: brom_out <= 64'd2151578802008365031;
    12'd463: brom_out <= 64'd3818591566592158579;
    12'd464: brom_out <= 64'd221168427156668620;
    12'd465: brom_out <= 64'd2432010159645715397;
    12'd466: brom_out <= 64'd7985210005529564458;
    12'd467: brom_out <= 64'd7521624398464494394;
    12'd468: brom_out <= 64'd6954602674252549157;
    12'd469: brom_out <= 64'd1772931732953384017;
    12'd470: brom_out <= 64'd3877069780779427166;
    12'd471: brom_out <= 64'd5821703083043290091;
    12'd472: brom_out <= 64'd5446263128435942946;
    12'd473: brom_out <= 64'd6209342773543205362;
    12'd474: brom_out <= 64'd8162841956676165738;
    12'd475: brom_out <= 64'd2739817607316069076;
    12'd476: brom_out <= 64'd5301890443195662787;
    12'd477: brom_out <= 64'd2802120147652768839;
    12'd478: brom_out <= 64'd1123132456013002459;
    12'd479: brom_out <= 64'd7701025136151381857;
    12'd480: brom_out <= 64'd3522401398456133729;
    12'd481: brom_out <= 64'd1121104267230146280;
    12'd482: brom_out <= 64'd4785516395754103712;
    12'd483: brom_out <= 64'd9204011995672087541;
    12'd484: brom_out <= 64'd6985849834050000541;
    12'd485: brom_out <= 64'd2806490387001446027;
    12'd486: brom_out <= 64'd6520183508896026597;
    12'd487: brom_out <= 64'd6903342917993908620;
    12'd488: brom_out <= 64'd7748187342122623094;
    12'd489: brom_out <= 64'd2145867268931626804;
    12'd490: brom_out <= 64'd6590112200699224071;
    12'd491: brom_out <= 64'd7207749336182051669;
    12'd492: brom_out <= 64'd4187235956733982846;
    12'd493: brom_out <= 64'd5209222732708414539;
    12'd494: brom_out <= 64'd4635191165656492150;
    12'd495: brom_out <= 64'd3079117042164723820;
    12'd496: brom_out <= 64'd9025502593406216690;
    12'd497: brom_out <= 64'd2137770580285350027;
    12'd498: brom_out <= 64'd5775523390321313615;
    12'd499: brom_out <= 64'd7086563346910060429;
    12'd500: brom_out <= 64'd1744638522500329828;
    12'd501: brom_out <= 64'd3442823001120628633;
    12'd502: brom_out <= 64'd3651945852037892795;
    12'd503: brom_out <= 64'd968497301989212927;
    12'd504: brom_out <= 64'd4533570374417505243;
    12'd505: brom_out <= 64'd5051377677337681721;
    12'd506: brom_out <= 64'd9097630694651455464;
    12'd507: brom_out <= 64'd2191685270051714447;
    12'd508: brom_out <= 64'd2914465977735506303;
    12'd509: brom_out <= 64'd5546600636589182767;
    12'd510: brom_out <= 64'd8074623464407446434;
    12'd511: brom_out <= 64'd8632183450091772719;
    12'd512: brom_out <= 64'd5976068779477487504;
    12'd513: brom_out <= 64'd4005117716490349010;
    12'd514: brom_out <= 64'd6744020006969895307;
    12'd515: brom_out <= 64'd5166836646587597065;
    12'd516: brom_out <= 64'd6061870125418198147;
    12'd517: brom_out <= 64'd1316412973703224049;
    12'd518: brom_out <= 64'd8927943298820454076;
    12'd519: brom_out <= 64'd6859486595377746448;
    12'd520: brom_out <= 64'd593042282816257658;
    12'd521: brom_out <= 64'd625448301026631026;
    12'd522: brom_out <= 64'd2799537887104471251;
    12'd523: brom_out <= 64'd6139871726171298472;
    12'd524: brom_out <= 64'd5181330732459777477;
    12'd525: brom_out <= 64'd5007472984365342136;
    12'd526: brom_out <= 64'd2187018093810691720;
    12'd527: brom_out <= 64'd6007025510947175156;
    12'd528: brom_out <= 64'd1271675644934090509;
    12'd529: brom_out <= 64'd2173064029340428803;
    12'd530: brom_out <= 64'd8522993162440537939;
    12'd531: brom_out <= 64'd2499747760317348668;
    12'd532: brom_out <= 64'd8013822734360034103;
    12'd533: brom_out <= 64'd666647422893437467;
    12'd534: brom_out <= 64'd5541375517500192895;
    12'd535: brom_out <= 64'd216156902476935823;
    12'd536: brom_out <= 64'd1177438167634269823;
    12'd537: brom_out <= 64'd2000665874345772028;
    12'd538: brom_out <= 64'd7698250944354989161;
    12'd539: brom_out <= 64'd516117442035369156;
    12'd540: brom_out <= 64'd6903674494547403458;
    12'd541: brom_out <= 64'd8577479475597382168;
    12'd542: brom_out <= 64'd5401614836719703272;
    12'd543: brom_out <= 64'd6143752504496732708;
    12'd544: brom_out <= 64'd8439932809411290039;
    12'd545: brom_out <= 64'd335350576825950082;
    12'd546: brom_out <= 64'd5152644225124011089;
    12'd547: brom_out <= 64'd7106724961015418341;
    12'd548: brom_out <= 64'd8791519766434938211;
    12'd549: brom_out <= 64'd6610019059717728193;
    12'd550: brom_out <= 64'd2868266086180312958;
    12'd551: brom_out <= 64'd7318335930499649148;
    12'd552: brom_out <= 64'd9170359323010223211;
    12'd553: brom_out <= 64'd7183671453211506471;
    12'd554: brom_out <= 64'd4765782474432323605;
    12'd555: brom_out <= 64'd6926826029504761109;
    12'd556: brom_out <= 64'd4794628727443279888;
    12'd557: brom_out <= 64'd3002431078669018093;
    12'd558: brom_out <= 64'd4633112736508198766;
    12'd559: brom_out <= 64'd5331734343637620507;
    12'd560: brom_out <= 64'd9036648888917473750;
    12'd561: brom_out <= 64'd4777872077056980363;
    12'd562: brom_out <= 64'd8336322066205089657;
    12'd563: brom_out <= 64'd6495472315871052654;
    12'd564: brom_out <= 64'd994064848121607400;
    12'd565: brom_out <= 64'd696331007242609412;
    12'd566: brom_out <= 64'd5410674334166473286;
    12'd567: brom_out <= 64'd6853549056042485036;
    12'd568: brom_out <= 64'd739218949392655402;
    12'd569: brom_out <= 64'd5951489724646106101;
    12'd570: brom_out <= 64'd8105253848644364450;
    12'd571: brom_out <= 64'd9087061851861541574;
    12'd572: brom_out <= 64'd7256022154194582960;
    12'd573: brom_out <= 64'd476664286229091365;
    12'd574: brom_out <= 64'd2464563482745670645;
    12'd575: brom_out <= 64'd6615395692181224670;
    12'd576: brom_out <= 64'd3874323780530106533;
    12'd577: brom_out <= 64'd1292420980917360603;
    12'd578: brom_out <= 64'd6351756831470743006;
    12'd579: brom_out <= 64'd7425855313841445797;
    12'd580: brom_out <= 64'd6928014622416298408;
    12'd581: brom_out <= 64'd7317450101610300559;
    12'd582: brom_out <= 64'd7747822092528642924;
    12'd583: brom_out <= 64'd8115948946013618884;
    12'd584: brom_out <= 64'd5718867093180509803;
    12'd585: brom_out <= 64'd3048930568431300260;
    12'd586: brom_out <= 64'd8252964877799973406;
    12'd587: brom_out <= 64'd3642980676160988416;
    12'd588: brom_out <= 64'd8433488676012520446;
    12'd589: brom_out <= 64'd8708749152152484117;
    12'd590: brom_out <= 64'd1481999355516963175;
    12'd591: brom_out <= 64'd1000681170679138810;
    12'd592: brom_out <= 64'd4363004334232094865;
    12'd593: brom_out <= 64'd8374712657994971746;
    12'd594: brom_out <= 64'd7137177962332868154;
    12'd595: brom_out <= 64'd5510182198338588319;
    12'd596: brom_out <= 64'd1021589499332145736;
    12'd597: brom_out <= 64'd7027237905526445895;
    12'd598: brom_out <= 64'd2857441601682776678;
    12'd599: brom_out <= 64'd3787408563903770001;
    12'd600: brom_out <= 64'd7929071200947786101;
    12'd601: brom_out <= 64'd2591362338410686344;
    12'd602: brom_out <= 64'd2703396381905810774;
    12'd603: brom_out <= 64'd9008273559910712642;
    12'd604: brom_out <= 64'd2663302601066611311;
    12'd605: brom_out <= 64'd6735328272190945037;
    12'd606: brom_out <= 64'd6034460869506398985;
    12'd607: brom_out <= 64'd3049253393215885299;
    12'd608: brom_out <= 64'd1085106348447748099;
    12'd609: brom_out <= 64'd6596423659328983517;
    12'd610: brom_out <= 64'd7280577718007746774;
    12'd611: brom_out <= 64'd4526467801563614800;
    12'd612: brom_out <= 64'd853076967703601242;
    12'd613: brom_out <= 64'd2788184500819922894;
    12'd614: brom_out <= 64'd8765870513679473211;
    12'd615: brom_out <= 64'd4057006210167085562;
    12'd616: brom_out <= 64'd809486194630696952;
    12'd617: brom_out <= 64'd9102526443833176819;
    12'd618: brom_out <= 64'd6768544696756439421;
    12'd619: brom_out <= 64'd5187244564822774566;
    12'd620: brom_out <= 64'd6179534021270744021;
    12'd621: brom_out <= 64'd4010273547781768614;
    12'd622: brom_out <= 64'd8658919390669651664;
    12'd623: brom_out <= 64'd8119863567815308140;
    12'd624: brom_out <= 64'd1403509903281381135;
    12'd625: brom_out <= 64'd5044057647806587586;
    12'd626: brom_out <= 64'd4551293125869120088;
    12'd627: brom_out <= 64'd8355797756938721784;
    12'd628: brom_out <= 64'd3510417462984237944;
    12'd629: brom_out <= 64'd5264632850253624255;
    12'd630: brom_out <= 64'd7524025148374291789;
    12'd631: brom_out <= 64'd1586452688103683977;
    12'd632: brom_out <= 64'd4619323584991910886;
    12'd633: brom_out <= 64'd2781981996128691817;
    12'd634: brom_out <= 64'd6326125611953081505;
    12'd635: brom_out <= 64'd5126919642324647453;
    12'd636: brom_out <= 64'd6415125647473131768;
    12'd637: brom_out <= 64'd3023184176706965674;
    12'd638: brom_out <= 64'd6658739335726264481;
    12'd639: brom_out <= 64'd5346911085079280798;
    12'd640: brom_out <= 64'd4066724171054462909;
    12'd641: brom_out <= 64'd3633979900330440892;
    12'd642: brom_out <= 64'd548261701981485419;
    12'd643: brom_out <= 64'd5832136871207562377;
    12'd644: brom_out <= 64'd1611893969776626643;
    12'd645: brom_out <= 64'd3822681420997167602;
    12'd646: brom_out <= 64'd9004572314107590138;
    12'd647: brom_out <= 64'd13846368282169064;
    12'd648: brom_out <= 64'd3603203538984367077;
    12'd649: brom_out <= 64'd1313331331708123806;
    12'd650: brom_out <= 64'd2805030511231525764;
    12'd651: brom_out <= 64'd585413331536420342;
    12'd652: brom_out <= 64'd8041554051968754776;
    12'd653: brom_out <= 64'd189106268087547237;
    12'd654: brom_out <= 64'd4806777613109574958;
    12'd655: brom_out <= 64'd1637309547778421810;
    12'd656: brom_out <= 64'd4710964611444245301;
    12'd657: brom_out <= 64'd7670512215868297688;
    12'd658: brom_out <= 64'd6926030477489072308;
    12'd659: brom_out <= 64'd1700990274694725704;
    12'd660: brom_out <= 64'd3118801396391702857;
    12'd661: brom_out <= 64'd3414624865495540060;
    12'd662: brom_out <= 64'd6265810223453665551;
    12'd663: brom_out <= 64'd4580895004721707237;
    12'd664: brom_out <= 64'd6828380608571071779;
    12'd665: brom_out <= 64'd3415602137400722566;
    12'd666: brom_out <= 64'd1512800906605612428;
    12'd667: brom_out <= 64'd581076090402175181;
    12'd668: brom_out <= 64'd8127637090793435339;
    12'd669: brom_out <= 64'd7025983680737965395;
    12'd670: brom_out <= 64'd4414284518212157732;
    12'd671: brom_out <= 64'd5129160045159717183;
    12'd672: brom_out <= 64'd8309796333647791448;
    12'd673: brom_out <= 64'd478119158814609466;
    12'd674: brom_out <= 64'd6457789071063052555;
    12'd675: brom_out <= 64'd9222684029687266857;
    12'd676: brom_out <= 64'd7940540358792163042;
    12'd677: brom_out <= 64'd2970910451624412054;
    12'd678: brom_out <= 64'd3823809497424801247;
    12'd679: brom_out <= 64'd8629179470676055812;
    12'd680: brom_out <= 64'd5684075750352032262;
    12'd681: brom_out <= 64'd7584921381365002484;
    12'd682: brom_out <= 64'd1415882188212200225;
    12'd683: brom_out <= 64'd5070366903226930676;
    12'd684: brom_out <= 64'd6468256505106281226;
    12'd685: brom_out <= 64'd5006322225260249573;
    12'd686: brom_out <= 64'd5300966512209250050;
    12'd687: brom_out <= 64'd1792685860936897610;
    12'd688: brom_out <= 64'd4441590473776765300;
    12'd689: brom_out <= 64'd7660349318066984762;
    12'd690: brom_out <= 64'd787340924847783803;
    12'd691: brom_out <= 64'd3544520116357534828;
    12'd692: brom_out <= 64'd8634381596625442610;
    12'd693: brom_out <= 64'd8020316467693061111;
    12'd694: brom_out <= 64'd7704688953664041795;
    12'd695: brom_out <= 64'd2993034213610705855;
    12'd696: brom_out <= 64'd6707938413484059878;
    12'd697: brom_out <= 64'd8250164011289223786;
    12'd698: brom_out <= 64'd1689924925158498949;
    12'd699: brom_out <= 64'd1418499548803264809;
    12'd700: brom_out <= 64'd8077069361822515059;
    12'd701: brom_out <= 64'd7935001385118833413;
    12'd702: brom_out <= 64'd6919778738676338510;
    12'd703: brom_out <= 64'd6867301955756113651;
    12'd704: brom_out <= 64'd2637886143940526168;
    12'd705: brom_out <= 64'd4912519834823704407;
    12'd706: brom_out <= 64'd7047875822701595031;
    12'd707: brom_out <= 64'd7129037378186886574;
    12'd708: brom_out <= 64'd4132551802894357262;
    12'd709: brom_out <= 64'd484472173182833754;
    12'd710: brom_out <= 64'd7687396513344217400;
    12'd711: brom_out <= 64'd6909328800562532699;
    12'd712: brom_out <= 64'd5320908759602881481;
    12'd713: brom_out <= 64'd2158981712364655228;
    12'd714: brom_out <= 64'd8135317976049821842;
    12'd715: brom_out <= 64'd2753317697438201979;
    12'd716: brom_out <= 64'd6222808144614635014;
    12'd717: brom_out <= 64'd760364662072605816;
    12'd718: brom_out <= 64'd5991839321352371775;
    12'd719: brom_out <= 64'd3039730646554404637;
    12'd720: brom_out <= 64'd7086452204833135780;
    12'd721: brom_out <= 64'd7605970516342646990;
    12'd722: brom_out <= 64'd1213734665504106333;
    12'd723: brom_out <= 64'd864420952012544153;
    12'd724: brom_out <= 64'd5695358218414993869;
    12'd725: brom_out <= 64'd1633105308011439896;
    12'd726: brom_out <= 64'd8240076708661524496;
    12'd727: brom_out <= 64'd1739832632716235247;
    12'd728: brom_out <= 64'd3372994486386929879;
    12'd729: brom_out <= 64'd6033457957159147088;
    12'd730: brom_out <= 64'd4519341334859734073;
    12'd731: brom_out <= 64'd1100322559612223103;
    12'd732: brom_out <= 64'd3022260544642597516;
    12'd733: brom_out <= 64'd1384350578725038654;
    12'd734: brom_out <= 64'd6353718731862795407;
    12'd735: brom_out <= 64'd2944315729599332973;
    12'd736: brom_out <= 64'd4291000205908552613;
    12'd737: brom_out <= 64'd3780203902726182378;
    12'd738: brom_out <= 64'd7224435870105783327;
    12'd739: brom_out <= 64'd6813168121181337925;
    12'd740: brom_out <= 64'd7819977419197775899;
    12'd741: brom_out <= 64'd984860808516397195;
    12'd742: brom_out <= 64'd7149484177775971227;
    12'd743: brom_out <= 64'd6230788417987498078;
    12'd744: brom_out <= 64'd1232654478032123658;
    12'd745: brom_out <= 64'd5375557945600039679;
    12'd746: brom_out <= 64'd196307236251518595;
    12'd747: brom_out <= 64'd6807433264447476885;
    12'd748: brom_out <= 64'd7099443897569798910;
    12'd749: brom_out <= 64'd4774005550677405386;
    12'd750: brom_out <= 64'd1364531386125093388;
    12'd751: brom_out <= 64'd4612786026804496290;
    12'd752: brom_out <= 64'd6665838607271236324;
    12'd753: brom_out <= 64'd9051064044881936071;
    12'd754: brom_out <= 64'd3633365094721677201;
    12'd755: brom_out <= 64'd6303308488427599573;
    12'd756: brom_out <= 64'd1297339388260599077;
    12'd757: brom_out <= 64'd1096701672734617714;
    12'd758: brom_out <= 64'd4041634879120597886;
    12'd759: brom_out <= 64'd4228600194548570995;
    12'd760: brom_out <= 64'd4070504440077246346;
    12'd761: brom_out <= 64'd2327416570468869961;
    12'd762: brom_out <= 64'd5917399405983790504;
    12'd763: brom_out <= 64'd8636091743291140867;
    12'd764: brom_out <= 64'd7603550242876584926;
    12'd765: brom_out <= 64'd6751843302554367241;
    12'd766: brom_out <= 64'd7094683365482870580;
    12'd767: brom_out <= 64'd1405441374437402737;
    12'd768: brom_out <= 64'd5792979130194094298;
    12'd769: brom_out <= 64'd78521125945926901;
    12'd770: brom_out <= 64'd1390063910113207289;
    12'd771: brom_out <= 64'd5823169037746669754;
    12'd772: brom_out <= 64'd4452291514428477137;
    12'd773: brom_out <= 64'd2984424569790546779;
    12'd774: brom_out <= 64'd7817367043308214467;
    12'd775: brom_out <= 64'd2826193018771081104;
    12'd776: brom_out <= 64'd222968537858942369;
    12'd777: brom_out <= 64'd402155676505531812;
    12'd778: brom_out <= 64'd1539629244627310107;
    12'd779: brom_out <= 64'd331508909586663393;
    12'd780: brom_out <= 64'd6650157038584548422;
    12'd781: brom_out <= 64'd2108314857132696248;
    12'd782: brom_out <= 64'd2456301622261705551;
    12'd783: brom_out <= 64'd4314974606150836240;
    12'd784: brom_out <= 64'd5318975219191802577;
    12'd785: brom_out <= 64'd25138778867551862;
    12'd786: brom_out <= 64'd8995741913985100290;
    12'd787: brom_out <= 64'd6191071447783597483;
    12'd788: brom_out <= 64'd4110541742333500737;
    12'd789: brom_out <= 64'd6925859408854431027;
    12'd790: brom_out <= 64'd7055503816228831091;
    12'd791: brom_out <= 64'd2851277803142913097;
    12'd792: brom_out <= 64'd5000944239179137954;
    12'd793: brom_out <= 64'd3941823019222225634;
    12'd794: brom_out <= 64'd5215707159989682948;
    12'd795: brom_out <= 64'd1649380730009983717;
    12'd796: brom_out <= 64'd1059548844895002697;
    12'd797: brom_out <= 64'd2104513439566953500;
    12'd798: brom_out <= 64'd5359119263554810248;
    12'd799: brom_out <= 64'd2937264643500724946;
    12'd800: brom_out <= 64'd5596038778869841895;
    12'd801: brom_out <= 64'd6162069774348355978;
    12'd802: brom_out <= 64'd1852954710699492504;
    12'd803: brom_out <= 64'd1088076550595330003;
    12'd804: brom_out <= 64'd7803653637595225642;
    12'd805: brom_out <= 64'd4039886054006184193;
    12'd806: brom_out <= 64'd4446551631123665655;
    12'd807: brom_out <= 64'd4530139836433554292;
    12'd808: brom_out <= 64'd3365288337767276247;
    12'd809: brom_out <= 64'd1368828974385072222;
    12'd810: brom_out <= 64'd6519885780090122409;
    12'd811: brom_out <= 64'd3515341576481069642;
    12'd812: brom_out <= 64'd5892854050328892876;
    12'd813: brom_out <= 64'd2548864131226053734;
    12'd814: brom_out <= 64'd2086211756656440867;
    12'd815: brom_out <= 64'd1191926010696125333;
    12'd816: brom_out <= 64'd6458351418566661432;
    12'd817: brom_out <= 64'd5693674981823269218;
    12'd818: brom_out <= 64'd2721341105491390085;
    12'd819: brom_out <= 64'd5447452542047891116;
    12'd820: brom_out <= 64'd4456208975303951299;
    12'd821: brom_out <= 64'd4023808547623250577;
    12'd822: brom_out <= 64'd5852786553912777685;
    12'd823: brom_out <= 64'd6096433046458680369;
    12'd824: brom_out <= 64'd5293457782313866956;
    12'd825: brom_out <= 64'd5860301030137744471;
    12'd826: brom_out <= 64'd1503390632805335282;
    12'd827: brom_out <= 64'd7516231720080428053;
    12'd828: brom_out <= 64'd2351375173829121150;
    12'd829: brom_out <= 64'd5598236424952292337;
    12'd830: brom_out <= 64'd8759164961417563512;
    12'd831: brom_out <= 64'd2099379525012808838;
    12'd832: brom_out <= 64'd2737158020017696281;
    12'd833: brom_out <= 64'd3950582044138852963;
    12'd834: brom_out <= 64'd6640287097552321424;
    12'd835: brom_out <= 64'd5402496919907892894;
    12'd836: brom_out <= 64'd2487979883454043411;
    12'd837: brom_out <= 64'd4977195593406246853;
    12'd838: brom_out <= 64'd17521832455993642;
    12'd839: brom_out <= 64'd1485900908579781315;
    12'd840: brom_out <= 64'd5607163649712091882;
    12'd841: brom_out <= 64'd7169512332837823604;
    12'd842: brom_out <= 64'd4217348036314092382;
    12'd843: brom_out <= 64'd5075818161597640077;
    12'd844: brom_out <= 64'd6229174968075775630;
    12'd845: brom_out <= 64'd3671551594854379962;
    12'd846: brom_out <= 64'd2051998054788366270;
    12'd847: brom_out <= 64'd2896324170644098685;
    12'd848: brom_out <= 64'd2216455649141208680;
    12'd849: brom_out <= 64'd4802317643994205088;
    12'd850: brom_out <= 64'd6796227057672368420;
    12'd851: brom_out <= 64'd8876448235781091709;
    12'd852: brom_out <= 64'd1314986123610772272;
    12'd853: brom_out <= 64'd1204415582446106112;
    12'd854: brom_out <= 64'd5880920423784685274;
    12'd855: brom_out <= 64'd6904517509735436689;
    12'd856: brom_out <= 64'd1455837426791755297;
    12'd857: brom_out <= 64'd830772712952438644;
    12'd858: brom_out <= 64'd6481798364871042424;
    12'd859: brom_out <= 64'd2634628254352179088;
    12'd860: brom_out <= 64'd1701272341948035267;
    12'd861: brom_out <= 64'd6640817230316013339;
    12'd862: brom_out <= 64'd1168596851321766456;
    12'd863: brom_out <= 64'd968559680937005248;
    12'd864: brom_out <= 64'd6071971305117248446;
    12'd865: brom_out <= 64'd8932324166801541824;
    12'd866: brom_out <= 64'd211205323560102598;
    12'd867: brom_out <= 64'd813325539083547321;
    12'd868: brom_out <= 64'd8108747189882628079;
    12'd869: brom_out <= 64'd326628130286763688;
    12'd870: brom_out <= 64'd962867634407305569;
    12'd871: brom_out <= 64'd1290930582866351128;
    12'd872: brom_out <= 64'd2023644405886518221;
    12'd873: brom_out <= 64'd1933497862117067950;
    12'd874: brom_out <= 64'd8948912045682648319;
    12'd875: brom_out <= 64'd5758110218168465728;
    12'd876: brom_out <= 64'd6396414439770314375;
    12'd877: brom_out <= 64'd8292868431172674679;
    12'd878: brom_out <= 64'd6259526245218962991;
    12'd879: brom_out <= 64'd1415788218295337537;
    12'd880: brom_out <= 64'd4050420130283138042;
    12'd881: brom_out <= 64'd5896964627131169131;
    12'd882: brom_out <= 64'd6160499120912117934;
    12'd883: brom_out <= 64'd2167999302398932480;
    12'd884: brom_out <= 64'd7977797132770592727;
    12'd885: brom_out <= 64'd6062567962812957720;
    12'd886: brom_out <= 64'd6552355050471698204;
    12'd887: brom_out <= 64'd3864165031077615023;
    12'd888: brom_out <= 64'd5243772136807645099;
    12'd889: brom_out <= 64'd7607391407196645499;
    12'd890: brom_out <= 64'd3651142297411659187;
    12'd891: brom_out <= 64'd6030263012495362676;
    12'd892: brom_out <= 64'd2314914454150418602;
    12'd893: brom_out <= 64'd4337748426843001873;
    12'd894: brom_out <= 64'd801305510105442737;
    12'd895: brom_out <= 64'd8460182789291736091;
    12'd896: brom_out <= 64'd2803267708398697040;
    12'd897: brom_out <= 64'd1514057220951852292;
    12'd898: brom_out <= 64'd4568079005623157455;
    12'd899: brom_out <= 64'd9117853174285888050;
    12'd900: brom_out <= 64'd8376944661285632772;
    12'd901: brom_out <= 64'd8804964526763484820;
    12'd902: brom_out <= 64'd8566281893646113;
    12'd903: brom_out <= 64'd3123787049644773702;
    12'd904: brom_out <= 64'd1618067356643750162;
    12'd905: brom_out <= 64'd502463928244531822;
    12'd906: brom_out <= 64'd3507173358449499779;
    12'd907: brom_out <= 64'd6797135268318975993;
    12'd908: brom_out <= 64'd2784388700362841711;
    12'd909: brom_out <= 64'd4101511390806188959;
    12'd910: brom_out <= 64'd6295273620685999449;
    12'd911: brom_out <= 64'd8303740360864384825;
    12'd912: brom_out <= 64'd4083878445077305523;
    12'd913: brom_out <= 64'd3183672025538269624;
    12'd914: brom_out <= 64'd2848313604941519881;
    12'd915: brom_out <= 64'd4648179036277464614;
    12'd916: brom_out <= 64'd6337223876791081151;
    12'd917: brom_out <= 64'd2699311646597186707;
    12'd918: brom_out <= 64'd7990560214861353583;
    12'd919: brom_out <= 64'd8130859604558591146;
    12'd920: brom_out <= 64'd7741923924364988008;
    12'd921: brom_out <= 64'd1673469281655632698;
    12'd922: brom_out <= 64'd1144176920185415535;
    12'd923: brom_out <= 64'd3249217722349422785;
    12'd924: brom_out <= 64'd2215604315896092670;
    12'd925: brom_out <= 64'd2714382757628886923;
    12'd926: brom_out <= 64'd2608525535082964773;
    12'd927: brom_out <= 64'd7657127696980843717;
    12'd928: brom_out <= 64'd3003943219615574075;
    12'd929: brom_out <= 64'd4024235301766674686;
    12'd930: brom_out <= 64'd47740789800497965;
    12'd931: brom_out <= 64'd4867650036211325578;
    12'd932: brom_out <= 64'd1382872280811698552;
    12'd933: brom_out <= 64'd2864923865331435467;
    12'd934: brom_out <= 64'd1901574174662490027;
    12'd935: brom_out <= 64'd9208255149800298927;
    12'd936: brom_out <= 64'd2803062370827609981;
    12'd937: brom_out <= 64'd8852578436638496032;
    12'd938: brom_out <= 64'd1992283337758212979;
    12'd939: brom_out <= 64'd2784125964689156344;
    12'd940: brom_out <= 64'd7700372050315114363;
    12'd941: brom_out <= 64'd1193634655463454607;
    12'd942: brom_out <= 64'd2875223919672073068;
    12'd943: brom_out <= 64'd4858729015412237653;
    12'd944: brom_out <= 64'd6019869478886392755;
    12'd945: brom_out <= 64'd1083320007172303764;
    12'd946: brom_out <= 64'd7140722186488696864;
    12'd947: brom_out <= 64'd456706321385894513;
    12'd948: brom_out <= 64'd6761610796267635122;
    12'd949: brom_out <= 64'd4372612876602253599;
    12'd950: brom_out <= 64'd3287964157657373940;
    12'd951: brom_out <= 64'd3815719428901871649;
    12'd952: brom_out <= 64'd5746142847633122703;
    12'd953: brom_out <= 64'd3617854177990257081;
    12'd954: brom_out <= 64'd3343459330700479572;
    12'd955: brom_out <= 64'd2333919523156828507;
    12'd956: brom_out <= 64'd3130462232530454679;
    12'd957: brom_out <= 64'd23757372729667867;
    12'd958: brom_out <= 64'd6889879677402930206;
    12'd959: brom_out <= 64'd3294907764858559824;
    12'd960: brom_out <= 64'd1065160304167154726;
    12'd961: brom_out <= 64'd7222535658536760892;
    12'd962: brom_out <= 64'd8625960684678229166;
    12'd963: brom_out <= 64'd8372383270641797411;
    12'd964: brom_out <= 64'd6953881865491377297;
    12'd965: brom_out <= 64'd2460547664794426212;
    12'd966: brom_out <= 64'd1707361404853655714;
    12'd967: brom_out <= 64'd8279003718731922783;
    12'd968: brom_out <= 64'd8151167855892330172;
    12'd969: brom_out <= 64'd4852120695248117336;
    12'd970: brom_out <= 64'd4633933436842356737;
    12'd971: brom_out <= 64'd587698803814343080;
    12'd972: brom_out <= 64'd4976637449741390052;
    12'd973: brom_out <= 64'd2544517863417907900;
    12'd974: brom_out <= 64'd6447223936141958870;
    12'd975: brom_out <= 64'd6219209598344493322;
    12'd976: brom_out <= 64'd3598379093835291182;
    12'd977: brom_out <= 64'd4082435061276421983;
    12'd978: brom_out <= 64'd3473787664538686576;
    12'd979: brom_out <= 64'd3440900081023092332;
    12'd980: brom_out <= 64'd3659981058207187100;
    12'd981: brom_out <= 64'd2264251713198501895;
    12'd982: brom_out <= 64'd8632467951852587989;
    12'd983: brom_out <= 64'd3154382174460298506;
    12'd984: brom_out <= 64'd4667723862850537194;
    12'd985: brom_out <= 64'd1179965516540825048;
    12'd986: brom_out <= 64'd3936667969893923919;
    12'd987: brom_out <= 64'd1704950911325584250;
    12'd988: brom_out <= 64'd9119962653750090131;
    12'd989: brom_out <= 64'd996377262630989551;
    12'd990: brom_out <= 64'd168302224660410828;
    12'd991: brom_out <= 64'd693939813520258859;
    12'd992: brom_out <= 64'd4910995540748981844;
    12'd993: brom_out <= 64'd4011863120442953560;
    12'd994: brom_out <= 64'd3657039766247532725;
    12'd995: brom_out <= 64'd5294995080171998451;
    12'd996: brom_out <= 64'd6432548891759686389;
    12'd997: brom_out <= 64'd6321448948253248513;
    12'd998: brom_out <= 64'd9123574294358671657;
    12'd999: brom_out <= 64'd3039518500019049569;
    12'd1000: brom_out <= 64'd9009408318896786413;
    12'd1001: brom_out <= 64'd6255317374299378826;
    12'd1002: brom_out <= 64'd3633265221550976288;
    12'd1003: brom_out <= 64'd7385984052681800207;
    12'd1004: brom_out <= 64'd5184317378868141180;
    12'd1005: brom_out <= 64'd592321105965206016;
    12'd1006: brom_out <= 64'd6244689180377020923;
    12'd1007: brom_out <= 64'd287410934104796108;
    12'd1008: brom_out <= 64'd8856063189815385885;
    12'd1009: brom_out <= 64'd6989967860725554358;
    12'd1010: brom_out <= 64'd1118592617708714057;
    12'd1011: brom_out <= 64'd5653837848356806718;
    12'd1012: brom_out <= 64'd5590202575696230393;
    12'd1013: brom_out <= 64'd3793296266665166283;
    12'd1014: brom_out <= 64'd3794573246885287845;
    12'd1015: brom_out <= 64'd6231911985272121732;
    12'd1016: brom_out <= 64'd4891968351182874667;
    12'd1017: brom_out <= 64'd6195679539347534888;
    12'd1018: brom_out <= 64'd8063678981840380015;
    12'd1019: brom_out <= 64'd4987501261148305465;
    12'd1020: brom_out <= 64'd5145477708918912727;
    12'd1021: brom_out <= 64'd792070567551351799;
    12'd1022: brom_out <= 64'd7920910159561005345;
    12'd1023: brom_out <= 64'd631785061731105457;
    12'd1024: brom_out <= 64'd6551015095526749063;
    12'd1025: brom_out <= 64'd4595731803495303327;
    12'd1026: brom_out <= 64'd8288530531944855590;
    12'd1027: brom_out <= 64'd3173670304377726411;
    12'd1028: brom_out <= 64'd8652315721870189437;
    12'd1029: brom_out <= 64'd1916386186435381995;
    12'd1030: brom_out <= 64'd6914660438246835908;
    12'd1031: brom_out <= 64'd4784390490314142871;
    12'd1032: brom_out <= 64'd3796382495133268725;
    12'd1033: brom_out <= 64'd1938270965119171169;
    12'd1034: brom_out <= 64'd2726913976235435110;
    12'd1035: brom_out <= 64'd7543858027698518528;
    12'd1036: brom_out <= 64'd15243861875148476;
    12'd1037: brom_out <= 64'd5349760899881279278;
    12'd1038: brom_out <= 64'd4148280298264435145;
    12'd1039: brom_out <= 64'd5390736926471664788;
    12'd1040: brom_out <= 64'd4040899244153570090;
    12'd1041: brom_out <= 64'd164674200546607604;
    12'd1042: brom_out <= 64'd4512365403662406081;
    12'd1043: brom_out <= 64'd6615260160847664585;
    12'd1044: brom_out <= 64'd2240211916433264831;
    12'd1045: brom_out <= 64'd6779561190491316855;
    12'd1046: brom_out <= 64'd7160540774931803866;
    12'd1047: brom_out <= 64'd6015795952029749156;
    12'd1048: brom_out <= 64'd5683041679221725246;
    12'd1049: brom_out <= 64'd8216051810600487589;
    12'd1050: brom_out <= 64'd9206702681534441482;
    12'd1051: brom_out <= 64'd5981994135735259692;
    12'd1052: brom_out <= 64'd8708624953667028585;
    12'd1053: brom_out <= 64'd8823402378843521219;
    12'd1054: brom_out <= 64'd7835211644950567469;
    12'd1055: brom_out <= 64'd5581925567248425011;
    12'd1056: brom_out <= 64'd284038871857826017;
    12'd1057: brom_out <= 64'd5218202542817394251;
    12'd1058: brom_out <= 64'd1445608483214028307;
    12'd1059: brom_out <= 64'd2520132840412007274;
    12'd1060: brom_out <= 64'd7096948766236504610;
    12'd1061: brom_out <= 64'd6050565049864378024;
    12'd1062: brom_out <= 64'd1778468342386166084;
    12'd1063: brom_out <= 64'd8104824511528610961;
    12'd1064: brom_out <= 64'd2554384204381077376;
    12'd1065: brom_out <= 64'd1556515623451888075;
    12'd1066: brom_out <= 64'd7537176118984402773;
    12'd1067: brom_out <= 64'd3261485979621056498;
    12'd1068: brom_out <= 64'd6463166748036722757;
    12'd1069: brom_out <= 64'd5548372674297715787;
    12'd1070: brom_out <= 64'd7664280676247221904;
    12'd1071: brom_out <= 64'd8163551390154089839;
    12'd1072: brom_out <= 64'd2529239563039080875;
    12'd1073: brom_out <= 64'd3161833067360455250;
    12'd1074: brom_out <= 64'd5407047594096528025;
    12'd1075: brom_out <= 64'd2122828736867373768;
    12'd1076: brom_out <= 64'd3847574256498121621;
    12'd1077: brom_out <= 64'd3248329190411644841;
    12'd1078: brom_out <= 64'd8373705960209865750;
    12'd1079: brom_out <= 64'd5096141494837811524;
    12'd1080: brom_out <= 64'd9106909176665937792;
    12'd1081: brom_out <= 64'd1021692220188325535;
    12'd1082: brom_out <= 64'd1100339483998246003;
    12'd1083: brom_out <= 64'd371088353612679558;
    12'd1084: brom_out <= 64'd111332146913263916;
    12'd1085: brom_out <= 64'd162862229894596551;
    12'd1086: brom_out <= 64'd849306692269551679;
    12'd1087: brom_out <= 64'd5417023988817079832;
    12'd1088: brom_out <= 64'd8872444489401680815;
    12'd1089: brom_out <= 64'd8400965878765427026;
    12'd1090: brom_out <= 64'd6943865764417683064;
    12'd1091: brom_out <= 64'd4082192015958411523;
    12'd1092: brom_out <= 64'd2343344652186686753;
    12'd1093: brom_out <= 64'd5351830350077338393;
    12'd1094: brom_out <= 64'd4751890286330071625;
    12'd1095: brom_out <= 64'd542606181224160151;
    12'd1096: brom_out <= 64'd4613289516563687559;
    12'd1097: brom_out <= 64'd2270794757509049429;
    12'd1098: brom_out <= 64'd806771516604876704;
    12'd1099: brom_out <= 64'd220166632239457975;
    12'd1100: brom_out <= 64'd6832924728641330482;
    12'd1101: brom_out <= 64'd8461937665451657542;
    12'd1102: brom_out <= 64'd6060747830154195747;
    12'd1103: brom_out <= 64'd6700911579012967260;
    12'd1104: brom_out <= 64'd2703826489472427745;
    12'd1105: brom_out <= 64'd5138973604269881666;
    12'd1106: brom_out <= 64'd3163609927867779470;
    12'd1107: brom_out <= 64'd8025602516218589744;
    12'd1108: brom_out <= 64'd3227682425404315158;
    12'd1109: brom_out <= 64'd259903952847149869;
    12'd1110: brom_out <= 64'd5069629123053312106;
    12'd1111: brom_out <= 64'd4014783758903962557;
    12'd1112: brom_out <= 64'd1952843272151728048;
    12'd1113: brom_out <= 64'd5800786890988034455;
    12'd1114: brom_out <= 64'd5757481406149589238;
    12'd1115: brom_out <= 64'd3414716947497933073;
    12'd1116: brom_out <= 64'd7104270022735541970;
    12'd1117: brom_out <= 64'd6105427606278424468;
    12'd1118: brom_out <= 64'd812235029203875617;
    12'd1119: brom_out <= 64'd7402170804642201058;
    12'd1120: brom_out <= 64'd2669547459691193432;
    12'd1121: brom_out <= 64'd6296175845735511856;
    12'd1122: brom_out <= 64'd1709606027938467824;
    12'd1123: brom_out <= 64'd4953097448697532735;
    12'd1124: brom_out <= 64'd4585039786213636068;
    12'd1125: brom_out <= 64'd1578854839664952686;
    12'd1126: brom_out <= 64'd5269356158780504864;
    12'd1127: brom_out <= 64'd198276819140143772;
    12'd1128: brom_out <= 64'd8345571030034495946;
    12'd1129: brom_out <= 64'd761655569867782735;
    12'd1130: brom_out <= 64'd5711684474143641757;
    12'd1131: brom_out <= 64'd9064173460967769874;
    12'd1132: brom_out <= 64'd6017550373169230213;
    12'd1133: brom_out <= 64'd7462540017383874819;
    12'd1134: brom_out <= 64'd8871767897380268353;
    12'd1135: brom_out <= 64'd7580464959537686266;
    12'd1136: brom_out <= 64'd538390155169630246;
    12'd1137: brom_out <= 64'd2206364998037189985;
    12'd1138: brom_out <= 64'd7452519829483945138;
    12'd1139: brom_out <= 64'd4812882446374196222;
    12'd1140: brom_out <= 64'd1458993785378647509;
    12'd1141: brom_out <= 64'd6548214732868127762;
    12'd1142: brom_out <= 64'd6524722060171723622;
    12'd1143: brom_out <= 64'd6200279617731237344;
    12'd1144: brom_out <= 64'd4078971191093288272;
    12'd1145: brom_out <= 64'd5584850174934109096;
    12'd1146: brom_out <= 64'd6501664496823873080;
    12'd1147: brom_out <= 64'd3805392669830113515;
    12'd1148: brom_out <= 64'd4583234557640069978;
    12'd1149: brom_out <= 64'd7110429745811052508;
    12'd1150: brom_out <= 64'd6382089802135409144;
    12'd1151: brom_out <= 64'd4463176173192127330;
    12'd1152: brom_out <= 64'd5908178380096272369;
    12'd1153: brom_out <= 64'd8061736108804448278;
    12'd1154: brom_out <= 64'd9103463721653978408;
    12'd1155: brom_out <= 64'd2822778535989408567;
    12'd1156: brom_out <= 64'd7993813175591520204;
    12'd1157: brom_out <= 64'd7721770747228916634;
    12'd1158: brom_out <= 64'd3032208211650146388;
    12'd1159: brom_out <= 64'd2295262262072788052;
    12'd1160: brom_out <= 64'd4682857295746554344;
    12'd1161: brom_out <= 64'd1873889101993027220;
    12'd1162: brom_out <= 64'd3139435852145256442;
    12'd1163: brom_out <= 64'd3457656149741362258;
    12'd1164: brom_out <= 64'd8934879803166669689;
    12'd1165: brom_out <= 64'd8744139465253655004;
    12'd1166: brom_out <= 64'd6846824846681755777;
    12'd1167: brom_out <= 64'd1606167506240542843;
    12'd1168: brom_out <= 64'd9076916340755116149;
    12'd1169: brom_out <= 64'd4886014524849036326;
    12'd1170: brom_out <= 64'd6610810496821611972;
    12'd1171: brom_out <= 64'd9032699219067860781;
    12'd1172: brom_out <= 64'd5024898852976039286;
    12'd1173: brom_out <= 64'd2403098808293565319;
    12'd1174: brom_out <= 64'd5041872014433074100;
    12'd1175: brom_out <= 64'd8647626436894153339;
    12'd1176: brom_out <= 64'd5040843640203270416;
    12'd1177: brom_out <= 64'd8869096447896116182;
    12'd1178: brom_out <= 64'd789422816571225780;
    12'd1179: brom_out <= 64'd3663232130631177082;
    12'd1180: brom_out <= 64'd4506204908127599502;
    12'd1181: brom_out <= 64'd6531604368224188806;
    12'd1182: brom_out <= 64'd4822808530417619233;
    12'd1183: brom_out <= 64'd8206033862314336179;
    12'd1184: brom_out <= 64'd1687335542159875606;
    12'd1185: brom_out <= 64'd8830493778383512291;
    12'd1186: brom_out <= 64'd9135823465542849361;
    12'd1187: brom_out <= 64'd2223491687363304360;
    12'd1188: brom_out <= 64'd6854317339658753350;
    12'd1189: brom_out <= 64'd4504726022688788972;
    12'd1190: brom_out <= 64'd7125835522680848670;
    12'd1191: brom_out <= 64'd9027321022514621789;
    12'd1192: brom_out <= 64'd8818463071528412136;
    12'd1193: brom_out <= 64'd2193863277718000910;
    12'd1194: brom_out <= 64'd5992435799082823388;
    12'd1195: brom_out <= 64'd6954783923074474543;
    12'd1196: brom_out <= 64'd7284478466022368184;
    12'd1197: brom_out <= 64'd5950625068259854648;
    12'd1198: brom_out <= 64'd176563187302484685;
    12'd1199: brom_out <= 64'd6714068005318992750;
    12'd1200: brom_out <= 64'd4938289008039594695;
    12'd1201: brom_out <= 64'd5258779288804072394;
    12'd1202: brom_out <= 64'd5802647509516054700;
    12'd1203: brom_out <= 64'd3642262225836421716;
    12'd1204: brom_out <= 64'd3688954750038363726;
    12'd1205: brom_out <= 64'd3885048787610312986;
    12'd1206: brom_out <= 64'd287090937624021185;
    12'd1207: brom_out <= 64'd7277929510343960039;
    12'd1208: brom_out <= 64'd6574977840107373503;
    12'd1209: brom_out <= 64'd1812932789727424157;
    12'd1210: brom_out <= 64'd7077564256689660660;
    12'd1211: brom_out <= 64'd8721513482441044300;
    12'd1212: brom_out <= 64'd821107918729627811;
    12'd1213: brom_out <= 64'd2520032607121689713;
    12'd1214: brom_out <= 64'd2749009972353655762;
    12'd1215: brom_out <= 64'd7804553392680594608;
    12'd1216: brom_out <= 64'd3547627594494878621;
    12'd1217: brom_out <= 64'd6265146028599173595;
    12'd1218: brom_out <= 64'd3136767173588347434;
    12'd1219: brom_out <= 64'd6250779680011007694;
    12'd1220: brom_out <= 64'd1549287551893278911;
    12'd1221: brom_out <= 64'd4675606206018073061;
    12'd1222: brom_out <= 64'd6579678929095156593;
    12'd1223: brom_out <= 64'd2052037289703534027;
    12'd1224: brom_out <= 64'd57560180524151836;
    12'd1225: brom_out <= 64'd3102877355736081607;
    12'd1226: brom_out <= 64'd8431525056773163324;
    12'd1227: brom_out <= 64'd5362137396733491930;
    12'd1228: brom_out <= 64'd7831437647304356508;
    12'd1229: brom_out <= 64'd4318098524395396650;
    12'd1230: brom_out <= 64'd25054386228368260;
    12'd1231: brom_out <= 64'd608396834745710365;
    12'd1232: brom_out <= 64'd5944864576936445287;
    12'd1233: brom_out <= 64'd3500901095250623076;
    12'd1234: brom_out <= 64'd978720527126678484;
    12'd1235: brom_out <= 64'd601771167641863668;
    12'd1236: brom_out <= 64'd5078991997579173257;
    12'd1237: brom_out <= 64'd1656312259292181257;
    12'd1238: brom_out <= 64'd5515184158531911546;
    12'd1239: brom_out <= 64'd8012349467558720615;
    12'd1240: brom_out <= 64'd684639643803771175;
    12'd1241: brom_out <= 64'd5084637108789426563;
    12'd1242: brom_out <= 64'd3281923340519708537;
    12'd1243: brom_out <= 64'd4722336290825604735;
    12'd1244: brom_out <= 64'd3340259218302706899;
    12'd1245: brom_out <= 64'd5700300283373190385;
    12'd1246: brom_out <= 64'd3591529433803820433;
    12'd1247: brom_out <= 64'd7912654433847146065;
    12'd1248: brom_out <= 64'd2468663283803736374;
    12'd1249: brom_out <= 64'd6205084145235084221;
    12'd1250: brom_out <= 64'd4585935009530136169;
    12'd1251: brom_out <= 64'd8880750789267131080;
    12'd1252: brom_out <= 64'd5798824876843371582;
    12'd1253: brom_out <= 64'd3516321696517407190;
    12'd1254: brom_out <= 64'd2212864360945965123;
    12'd1255: brom_out <= 64'd3975183427385598615;
    12'd1256: brom_out <= 64'd1837680713908133646;
    12'd1257: brom_out <= 64'd8931667155076678830;
    12'd1258: brom_out <= 64'd672919549451933827;
    12'd1259: brom_out <= 64'd7789650034503307067;
    12'd1260: brom_out <= 64'd2036591841189774695;
    12'd1261: brom_out <= 64'd5342489680170388343;
    12'd1262: brom_out <= 64'd6072046178105556475;
    12'd1263: brom_out <= 64'd2905515105513391987;
    12'd1264: brom_out <= 64'd1178188298187125443;
    12'd1265: brom_out <= 64'd5549144129026746013;
    12'd1266: brom_out <= 64'd5545686084666219710;
    12'd1267: brom_out <= 64'd1343223045376093288;
    12'd1268: brom_out <= 64'd3110559949174149380;
    12'd1269: brom_out <= 64'd3733261563727931026;
    12'd1270: brom_out <= 64'd1330381704714286085;
    12'd1271: brom_out <= 64'd36022640168924989;
    12'd1272: brom_out <= 64'd5873106135293020355;
    12'd1273: brom_out <= 64'd4076427909784645200;
    12'd1274: brom_out <= 64'd1435120993511282705;
    12'd1275: brom_out <= 64'd995086951603849713;
    12'd1276: brom_out <= 64'd8803778985884906727;
    12'd1277: brom_out <= 64'd4287893524448971608;
    12'd1278: brom_out <= 64'd6585546512385483974;
    12'd1279: brom_out <= 64'd5602381032211604622;
    12'd1280: brom_out <= 64'd2991444385089030097;
    12'd1281: brom_out <= 64'd3256237472906815544;
    12'd1282: brom_out <= 64'd6427097281726706628;
    12'd1283: brom_out <= 64'd4184126388409380134;
    12'd1284: brom_out <= 64'd4183299227927339195;
    12'd1285: brom_out <= 64'd3895031829224767346;
    12'd1286: brom_out <= 64'd3119079411128405209;
    12'd1287: brom_out <= 64'd9155661255527747178;
    12'd1288: brom_out <= 64'd1122397655549924356;
    12'd1289: brom_out <= 64'd2310560732345386485;
    12'd1290: brom_out <= 64'd5564951036314476973;
    12'd1291: brom_out <= 64'd7216537363218896285;
    12'd1292: brom_out <= 64'd2527297775950676908;
    12'd1293: brom_out <= 64'd634583883983266145;
    12'd1294: brom_out <= 64'd3036875632463858834;
    12'd1295: brom_out <= 64'd2242810203672903028;
    12'd1296: brom_out <= 64'd6281663284576107517;
    12'd1297: brom_out <= 64'd8897863336940776164;
    12'd1298: brom_out <= 64'd4794722994419500598;
    12'd1299: brom_out <= 64'd6643848106357390455;
    12'd1300: brom_out <= 64'd7533491753178725717;
    12'd1301: brom_out <= 64'd8963917332809987708;
    12'd1302: brom_out <= 64'd8580562440646539131;
    12'd1303: brom_out <= 64'd3047197073143512046;
    12'd1304: brom_out <= 64'd8697599446790123293;
    12'd1305: brom_out <= 64'd7216151128053990306;
    12'd1306: brom_out <= 64'd5318448438505440257;
    12'd1307: brom_out <= 64'd1341898580837423017;
    12'd1308: brom_out <= 64'd235142833563334451;
    12'd1309: brom_out <= 64'd8903487350221356454;
    12'd1310: brom_out <= 64'd1078913570171309648;
    12'd1311: brom_out <= 64'd8356640971005957295;
    12'd1312: brom_out <= 64'd8124953238658307565;
    12'd1313: brom_out <= 64'd4346661030238530214;
    12'd1314: brom_out <= 64'd6514515671117556603;
    12'd1315: brom_out <= 64'd1393076932459315047;
    12'd1316: brom_out <= 64'd5808776274764837854;
    12'd1317: brom_out <= 64'd5245797325928432520;
    12'd1318: brom_out <= 64'd1737665055851572803;
    12'd1319: brom_out <= 64'd2418821237100432937;
    12'd1320: brom_out <= 64'd4625294087119433729;
    12'd1321: brom_out <= 64'd593907935894979160;
    12'd1322: brom_out <= 64'd3148801124557623449;
    12'd1323: brom_out <= 64'd4335064197964659539;
    12'd1324: brom_out <= 64'd75966845172534173;
    12'd1325: brom_out <= 64'd1400719953817300295;
    12'd1326: brom_out <= 64'd1113248537812598346;
    12'd1327: brom_out <= 64'd6536107692361147554;
    12'd1328: brom_out <= 64'd5782598045554155253;
    12'd1329: brom_out <= 64'd8155382693858119578;
    12'd1330: brom_out <= 64'd1141036854004408858;
    12'd1331: brom_out <= 64'd4889370594359438957;
    12'd1332: brom_out <= 64'd7870108581299121483;
    12'd1333: brom_out <= 64'd6814376656091464033;
    12'd1334: brom_out <= 64'd4196968460687196785;
    12'd1335: brom_out <= 64'd7707838255361434376;
    12'd1336: brom_out <= 64'd5991059833680697521;
    12'd1337: brom_out <= 64'd5811578762429694397;
    12'd1338: brom_out <= 64'd4613903798598080436;
    12'd1339: brom_out <= 64'd1091320823777447142;
    12'd1340: brom_out <= 64'd8100294372597586432;
    12'd1341: brom_out <= 64'd2958152679937921299;
    12'd1342: brom_out <= 64'd3504473931275065124;
    12'd1343: brom_out <= 64'd4756412739101574244;
    12'd1344: brom_out <= 64'd9166670786663116443;
    12'd1345: brom_out <= 64'd8058518244289887562;
    12'd1346: brom_out <= 64'd5395617652967469222;
    12'd1347: brom_out <= 64'd5165561524482769986;
    12'd1348: brom_out <= 64'd7083423175763586691;
    12'd1349: brom_out <= 64'd2432890573058181033;
    12'd1350: brom_out <= 64'd7441158198174016671;
    12'd1351: brom_out <= 64'd4040582382191874932;
    12'd1352: brom_out <= 64'd7173654840489607776;
    12'd1353: brom_out <= 64'd7417372571204481830;
    12'd1354: brom_out <= 64'd8838718518559474163;
    12'd1355: brom_out <= 64'd5201503226485455237;
    12'd1356: brom_out <= 64'd1947243181919420491;
    12'd1357: brom_out <= 64'd8177505488046858016;
    12'd1358: brom_out <= 64'd3854484312171404456;
    12'd1359: brom_out <= 64'd2919958029833209633;
    12'd1360: brom_out <= 64'd3115848091286679823;
    12'd1361: brom_out <= 64'd7011739122720262005;
    12'd1362: brom_out <= 64'd8317588540207922448;
    12'd1363: brom_out <= 64'd2855397955646245100;
    12'd1364: brom_out <= 64'd5226535173943436928;
    12'd1365: brom_out <= 64'd8942074700439913039;
    12'd1366: brom_out <= 64'd3682273990606439039;
    12'd1367: brom_out <= 64'd7528195295407567929;
    12'd1368: brom_out <= 64'd750361034814781007;
    12'd1369: brom_out <= 64'd6146999979043876520;
    12'd1370: brom_out <= 64'd4397702267799328608;
    12'd1371: brom_out <= 64'd9000490380987386148;
    12'd1372: brom_out <= 64'd3592198641247208794;
    12'd1373: brom_out <= 64'd1425902537865729979;
    12'd1374: brom_out <= 64'd3433509905416311683;
    12'd1375: brom_out <= 64'd5471432485527519578;
    12'd1376: brom_out <= 64'd5654726277541044038;
    12'd1377: brom_out <= 64'd3512444620723338488;
    12'd1378: brom_out <= 64'd5083175541303528685;
    12'd1379: brom_out <= 64'd6738164926973299742;
    12'd1380: brom_out <= 64'd4510264232516592952;
    12'd1381: brom_out <= 64'd8955222256909707638;
    12'd1382: brom_out <= 64'd2931018764400806070;
    12'd1383: brom_out <= 64'd6888711580551652825;
    12'd1384: brom_out <= 64'd5208814341045079371;
    12'd1385: brom_out <= 64'd3962315922150850049;
    12'd1386: brom_out <= 64'd8312556079981528030;
    12'd1387: brom_out <= 64'd2509718512183293069;
    12'd1388: brom_out <= 64'd5551115908770807940;
    12'd1389: brom_out <= 64'd8052177048263815731;
    12'd1390: brom_out <= 64'd585096259269936048;
    12'd1391: brom_out <= 64'd6044746018222371047;
    12'd1392: brom_out <= 64'd3558399091024426444;
    12'd1393: brom_out <= 64'd962407481846958591;
    12'd1394: brom_out <= 64'd4322711149969805068;
    12'd1395: brom_out <= 64'd8140874147456852453;
    12'd1396: brom_out <= 64'd1491544262489362891;
    12'd1397: brom_out <= 64'd4231499661440202131;
    12'd1398: brom_out <= 64'd6079977503648451335;
    12'd1399: brom_out <= 64'd2450795518335383150;
    12'd1400: brom_out <= 64'd4764036910647300995;
    12'd1401: brom_out <= 64'd2686589714625351870;
    12'd1402: brom_out <= 64'd1985994961055839280;
    12'd1403: brom_out <= 64'd1882086957153388148;
    12'd1404: brom_out <= 64'd9197868711120196895;
    12'd1405: brom_out <= 64'd6524547434638763383;
    12'd1406: brom_out <= 64'd6769971139694742693;
    12'd1407: brom_out <= 64'd448403919027889030;
    12'd1408: brom_out <= 64'd7646914504675205489;
    12'd1409: brom_out <= 64'd8816500119098547526;
    12'd1410: brom_out <= 64'd8256294627998732981;
    12'd1411: brom_out <= 64'd563696475519026428;
    12'd1412: brom_out <= 64'd5713577346046003020;
    12'd1413: brom_out <= 64'd6458810129696068279;
    12'd1414: brom_out <= 64'd1478979661686592040;
    12'd1415: brom_out <= 64'd3489052947642352681;
    12'd1416: brom_out <= 64'd3065938557921374089;
    12'd1417: brom_out <= 64'd6566502495667702930;
    12'd1418: brom_out <= 64'd2610367100111832212;
    12'd1419: brom_out <= 64'd8878323482694811936;
    12'd1420: brom_out <= 64'd2744296939060575530;
    12'd1421: brom_out <= 64'd5790249722416355499;
    12'd1422: brom_out <= 64'd3368411057424669635;
    12'd1423: brom_out <= 64'd3703586401268449278;
    12'd1424: brom_out <= 64'd1555308162728177297;
    12'd1425: brom_out <= 64'd9161163982018377625;
    12'd1426: brom_out <= 64'd4054013996166535507;
    12'd1427: brom_out <= 64'd5562682736650988466;
    12'd1428: brom_out <= 64'd220088159844794260;
    12'd1429: brom_out <= 64'd539332076438600639;
    12'd1430: brom_out <= 64'd7976876523254192230;
    12'd1431: brom_out <= 64'd6277239556914161008;
    12'd1432: brom_out <= 64'd6550225160897858344;
    12'd1433: brom_out <= 64'd8513875384724119180;
    12'd1434: brom_out <= 64'd7892653319965062638;
    12'd1435: brom_out <= 64'd1584884239282854430;
    12'd1436: brom_out <= 64'd5490294517849368108;
    12'd1437: brom_out <= 64'd9079580109520213237;
    12'd1438: brom_out <= 64'd6199672516180526071;
    12'd1439: brom_out <= 64'd281616783970276541;
    12'd1440: brom_out <= 64'd2141707773911427712;
    12'd1441: brom_out <= 64'd3763494781935998767;
    12'd1442: brom_out <= 64'd635855831193566106;
    12'd1443: brom_out <= 64'd5253324035467520156;
    12'd1444: brom_out <= 64'd7593220218804307867;
    12'd1445: brom_out <= 64'd7207426732065879308;
    12'd1446: brom_out <= 64'd8341925111666110475;
    12'd1447: brom_out <= 64'd1472757774526024785;
    12'd1448: brom_out <= 64'd5418439566171715291;
    12'd1449: brom_out <= 64'd7445483466275733942;
    12'd1450: brom_out <= 64'd8673620925411977753;
    12'd1451: brom_out <= 64'd4594800911237165801;
    12'd1452: brom_out <= 64'd4249431574386262900;
    12'd1453: brom_out <= 64'd6403028868537790655;
    12'd1454: brom_out <= 64'd2847404267546166357;
    12'd1455: brom_out <= 64'd1519567052495348237;
    12'd1456: brom_out <= 64'd7010796944267998638;
    12'd1457: brom_out <= 64'd1314283965644365680;
    12'd1458: brom_out <= 64'd3468411571066471426;
    12'd1459: brom_out <= 64'd468569663261293589;
    12'd1460: brom_out <= 64'd7135696680823117604;
    12'd1461: brom_out <= 64'd2991053525981376065;
    12'd1462: brom_out <= 64'd6230035500739914156;
    12'd1463: brom_out <= 64'd4841250990366375746;
    12'd1464: brom_out <= 64'd8692551628537520016;
    12'd1465: brom_out <= 64'd132458694871421557;
    12'd1466: brom_out <= 64'd8513076200388136183;
    12'd1467: brom_out <= 64'd917141149160099628;
    12'd1468: brom_out <= 64'd4824069180043442917;
    12'd1469: brom_out <= 64'd8501478292815056322;
    12'd1470: brom_out <= 64'd1141842582310077908;
    12'd1471: brom_out <= 64'd3314498144052701739;
    12'd1472: brom_out <= 64'd4393262027419573708;
    12'd1473: brom_out <= 64'd6333478367606839407;
    12'd1474: brom_out <= 64'd3058650903359729066;
    12'd1475: brom_out <= 64'd7178172838362117853;
    12'd1476: brom_out <= 64'd8893614490103508778;
    12'd1477: brom_out <= 64'd671685460762616247;
    12'd1478: brom_out <= 64'd7462328687096900295;
    12'd1479: brom_out <= 64'd3897349523513245448;
    12'd1480: brom_out <= 64'd4159689793066360690;
    12'd1481: brom_out <= 64'd623780653727302203;
    12'd1482: brom_out <= 64'd6283534932199547339;
    12'd1483: brom_out <= 64'd8163830362846381072;
    12'd1484: brom_out <= 64'd654752926994167022;
    12'd1485: brom_out <= 64'd268999905903068517;
    12'd1486: brom_out <= 64'd6628447066861725489;
    12'd1487: brom_out <= 64'd2439176352400363216;
    12'd1488: brom_out <= 64'd4919595983980879989;
    12'd1489: brom_out <= 64'd7692433165927744565;
    12'd1490: brom_out <= 64'd6301640391988730655;
    12'd1491: brom_out <= 64'd8199554349178138502;
    12'd1492: brom_out <= 64'd2816403948006974041;
    12'd1493: brom_out <= 64'd5867286401481316597;
    12'd1494: brom_out <= 64'd8969075915070151768;
    12'd1495: brom_out <= 64'd3137606336581079208;
    12'd1496: brom_out <= 64'd4919750730687193807;
    12'd1497: brom_out <= 64'd7005569702398285466;
    12'd1498: brom_out <= 64'd8694371873892844208;
    12'd1499: brom_out <= 64'd8317491426765841036;
    12'd1500: brom_out <= 64'd4413826527383477878;
    12'd1501: brom_out <= 64'd6767449512620135517;
    12'd1502: brom_out <= 64'd7030554445186196665;
    12'd1503: brom_out <= 64'd3167893952487493944;
    12'd1504: brom_out <= 64'd5729951333194461427;
    12'd1505: brom_out <= 64'd1885864751055057353;
    12'd1506: brom_out <= 64'd7978110531043641769;
    12'd1507: brom_out <= 64'd9081318113255327118;
    12'd1508: brom_out <= 64'd8743332571195579934;
    12'd1509: brom_out <= 64'd2477351137960909314;
    12'd1510: brom_out <= 64'd9129774312610320619;
    12'd1511: brom_out <= 64'd6552917894363667778;
    12'd1512: brom_out <= 64'd2240289491309476277;
    12'd1513: brom_out <= 64'd426035889455316640;
    12'd1514: brom_out <= 64'd8440836487301065001;
    12'd1515: brom_out <= 64'd1389138119124998720;
    12'd1516: brom_out <= 64'd2173356542276770935;
    12'd1517: brom_out <= 64'd2013262658437665285;
    12'd1518: brom_out <= 64'd1755068967933061315;
    12'd1519: brom_out <= 64'd1885157749448756501;
    12'd1520: brom_out <= 64'd1376701315345052441;
    12'd1521: brom_out <= 64'd3707251717625885791;
    12'd1522: brom_out <= 64'd6593921752856366535;
    12'd1523: brom_out <= 64'd7071548278656136848;
    12'd1524: brom_out <= 64'd3167756150689666531;
    12'd1525: brom_out <= 64'd855970050860984344;
    12'd1526: brom_out <= 64'd3784018163499518601;
    12'd1527: brom_out <= 64'd8516443880759784307;
    12'd1528: brom_out <= 64'd5939667306004532036;
    12'd1529: brom_out <= 64'd1509886436569520070;
    12'd1530: brom_out <= 64'd7427050020511569441;
    12'd1531: brom_out <= 64'd2656374355877288154;
    12'd1532: brom_out <= 64'd2935114005611711057;
    12'd1533: brom_out <= 64'd6810071412848208525;
    12'd1534: brom_out <= 64'd7692930341342185952;
    12'd1535: brom_out <= 64'd6055970653617461320;
    12'd1536: brom_out <= 64'd3392617565049336557;
    12'd1537: brom_out <= 64'd2678065129254935256;
    12'd1538: brom_out <= 64'd7131970059357333029;
    12'd1539: brom_out <= 64'd1676519968667390242;
    12'd1540: brom_out <= 64'd2230049327513614869;
    12'd1541: brom_out <= 64'd4586326237824140186;
    12'd1542: brom_out <= 64'd3854526127297200834;
    12'd1543: brom_out <= 64'd6026366267866628186;
    12'd1544: brom_out <= 64'd7479147464852913991;
    12'd1545: brom_out <= 64'd2164118330631263854;
    12'd1546: brom_out <= 64'd5742128143480654282;
    12'd1547: brom_out <= 64'd4007459461997400903;
    12'd1548: brom_out <= 64'd7538107808473199530;
    12'd1549: brom_out <= 64'd5823730381839252049;
    12'd1550: brom_out <= 64'd822715829145346347;
    12'd1551: brom_out <= 64'd642913437998720848;
    12'd1552: brom_out <= 64'd2263269548655216762;
    12'd1553: brom_out <= 64'd7922160522628872772;
    12'd1554: brom_out <= 64'd3329822700088162495;
    12'd1555: brom_out <= 64'd220774408946330784;
    12'd1556: brom_out <= 64'd6798664954031634633;
    12'd1557: brom_out <= 64'd5058062501522262208;
    12'd1558: brom_out <= 64'd4175560118002252921;
    12'd1559: brom_out <= 64'd3173784488041209200;
    12'd1560: brom_out <= 64'd6982695801609760735;
    12'd1561: brom_out <= 64'd6798974422792108364;
    12'd1562: brom_out <= 64'd6913663135607926584;
    12'd1563: brom_out <= 64'd4700118327586250533;
    12'd1564: brom_out <= 64'd6068442745462420874;
    12'd1565: brom_out <= 64'd7122058084065222170;
    12'd1566: brom_out <= 64'd2228552985412019277;
    12'd1567: brom_out <= 64'd8078411340332537200;
    12'd1568: brom_out <= 64'd8216761589456164;
    12'd1569: brom_out <= 64'd3388698090164268880;
    12'd1570: brom_out <= 64'd5266018003312504579;
    12'd1571: brom_out <= 64'd1292270614421363347;
    12'd1572: brom_out <= 64'd9102413699342598757;
    12'd1573: brom_out <= 64'd8954948950927174815;
    12'd1574: brom_out <= 64'd3580819943894297764;
    12'd1575: brom_out <= 64'd3288117840036850138;
    12'd1576: brom_out <= 64'd6925371594294004533;
    12'd1577: brom_out <= 64'd5028445509124063333;
    12'd1578: brom_out <= 64'd4784055077466289542;
    12'd1579: brom_out <= 64'd6012239089180365601;
    12'd1580: brom_out <= 64'd1568136098664689522;
    12'd1581: brom_out <= 64'd8614484543584024473;
    12'd1582: brom_out <= 64'd4419790281338715805;
    12'd1583: brom_out <= 64'd4583713786487905006;
    12'd1584: brom_out <= 64'd8186964208105355814;
    12'd1585: brom_out <= 64'd5322751941608048097;
    12'd1586: brom_out <= 64'd8817464271798224027;
    12'd1587: brom_out <= 64'd615834550689196678;
    12'd1588: brom_out <= 64'd1676869911627098617;
    12'd1589: brom_out <= 64'd6235368745691702325;
    12'd1590: brom_out <= 64'd4401819749409430491;
    12'd1591: brom_out <= 64'd5204306756936923712;
    12'd1592: brom_out <= 64'd6849437044168275747;
    12'd1593: brom_out <= 64'd9036507672267599775;
    12'd1594: brom_out <= 64'd7286314464983170863;
    12'd1595: brom_out <= 64'd6118620384573872227;
    12'd1596: brom_out <= 64'd8444867741212273661;
    12'd1597: brom_out <= 64'd6729280471890946438;
    12'd1598: brom_out <= 64'd9151515973652221402;
    12'd1599: brom_out <= 64'd8810587607558976549;
    12'd1600: brom_out <= 64'd5039744181953194803;
    12'd1601: brom_out <= 64'd5959304096792569751;
    12'd1602: brom_out <= 64'd637799399688374479;
    12'd1603: brom_out <= 64'd1809521424258670838;
    12'd1604: brom_out <= 64'd3468732936118861906;
    12'd1605: brom_out <= 64'd6078180130894032113;
    12'd1606: brom_out <= 64'd2777986735042830839;
    12'd1607: brom_out <= 64'd2522336249437108104;
    12'd1608: brom_out <= 64'd3064309850488305304;
    12'd1609: brom_out <= 64'd716419806412526384;
    12'd1610: brom_out <= 64'd4131185556170130308;
    12'd1611: brom_out <= 64'd5182512363142578659;
    12'd1612: brom_out <= 64'd391518006782257654;
    12'd1613: brom_out <= 64'd3873551248534087511;
    12'd1614: brom_out <= 64'd2051836413390839457;
    12'd1615: brom_out <= 64'd2321442173369150588;
    12'd1616: brom_out <= 64'd5471972468712594632;
    12'd1617: brom_out <= 64'd6515807241519471828;
    12'd1618: brom_out <= 64'd8595678383967341286;
    12'd1619: brom_out <= 64'd7251072921457186698;
    12'd1620: brom_out <= 64'd8395167631823199941;
    12'd1621: brom_out <= 64'd2268799027509688551;
    12'd1622: brom_out <= 64'd8907923421314590115;
    12'd1623: brom_out <= 64'd6380806961761902536;
    12'd1624: brom_out <= 64'd6626178562688381462;
    12'd1625: brom_out <= 64'd6693195915515107207;
    12'd1626: brom_out <= 64'd5769552562384596599;
    12'd1627: brom_out <= 64'd6757311289111676977;
    12'd1628: brom_out <= 64'd9209536114756024834;
    12'd1629: brom_out <= 64'd3816207022314241251;
    12'd1630: brom_out <= 64'd8947667063148711049;
    12'd1631: brom_out <= 64'd1572212746857595784;
    12'd1632: brom_out <= 64'd1628906345678539120;
    12'd1633: brom_out <= 64'd9099378341091656482;
    12'd1634: brom_out <= 64'd1544674224130596118;
    12'd1635: brom_out <= 64'd704204137755443298;
    12'd1636: brom_out <= 64'd4368700210148671551;
    12'd1637: brom_out <= 64'd4997739833658486655;
    12'd1638: brom_out <= 64'd6319435406754674390;
    12'd1639: brom_out <= 64'd8315450962467588491;
    12'd1640: brom_out <= 64'd7705829573832500897;
    12'd1641: brom_out <= 64'd9178637669322844693;
    12'd1642: brom_out <= 64'd4677673593772524828;
    12'd1643: brom_out <= 64'd5227644328066207813;
    12'd1644: brom_out <= 64'd4934228471949137670;
    12'd1645: brom_out <= 64'd3024775562432476191;
    12'd1646: brom_out <= 64'd5511461520034253554;
    12'd1647: brom_out <= 64'd7613867444966436683;
    12'd1648: brom_out <= 64'd3528090222809025860;
    12'd1649: brom_out <= 64'd1745036897308546683;
    12'd1650: brom_out <= 64'd1607600945152906512;
    12'd1651: brom_out <= 64'd7080205292498256390;
    12'd1652: brom_out <= 64'd1258669831230654444;
    12'd1653: brom_out <= 64'd8687882850748879926;
    12'd1654: brom_out <= 64'd2170069437537526133;
    12'd1655: brom_out <= 64'd597184167161759606;
    12'd1656: brom_out <= 64'd8798316185508471405;
    12'd1657: brom_out <= 64'd3186873110017313996;
    12'd1658: brom_out <= 64'd7183585907134239486;
    12'd1659: brom_out <= 64'd1714483633892986712;
    12'd1660: brom_out <= 64'd6154077313509807261;
    12'd1661: brom_out <= 64'd8700108686837974136;
    12'd1662: brom_out <= 64'd4955822627172985255;
    12'd1663: brom_out <= 64'd3850279675568096104;
    12'd1664: brom_out <= 64'd1002059954001900696;
    12'd1665: brom_out <= 64'd4114200839665517402;
    12'd1666: brom_out <= 64'd4687421323741025393;
    12'd1667: brom_out <= 64'd3433750853083519277;
    12'd1668: brom_out <= 64'd2757773614559033666;
    12'd1669: brom_out <= 64'd3887545247412752285;
    12'd1670: brom_out <= 64'd4725094368207763061;
    12'd1671: brom_out <= 64'd270433545850009328;
    12'd1672: brom_out <= 64'd1490887556607246244;
    12'd1673: brom_out <= 64'd5792180516837140858;
    12'd1674: brom_out <= 64'd91987351604627050;
    12'd1675: brom_out <= 64'd7166490740407512639;
    12'd1676: brom_out <= 64'd7104811893195087792;
    12'd1677: brom_out <= 64'd5679738671843934604;
    12'd1678: brom_out <= 64'd7767226473893413332;
    12'd1679: brom_out <= 64'd4307950442227902464;
    12'd1680: brom_out <= 64'd307156682351195017;
    12'd1681: brom_out <= 64'd3393684384123953368;
    12'd1682: brom_out <= 64'd4898893176619253892;
    12'd1683: brom_out <= 64'd4572460370399290474;
    12'd1684: brom_out <= 64'd8730278730941939396;
    12'd1685: brom_out <= 64'd5238391540599559172;
    12'd1686: brom_out <= 64'd3005741243809146285;
    12'd1687: brom_out <= 64'd5586233649254080813;
    12'd1688: brom_out <= 64'd3107918471259441615;
    12'd1689: brom_out <= 64'd585382463249167719;
    12'd1690: brom_out <= 64'd725251043603134492;
    12'd1691: brom_out <= 64'd2221481776280657367;
    12'd1692: brom_out <= 64'd6460685242337216620;
    12'd1693: brom_out <= 64'd62214353023950165;
    12'd1694: brom_out <= 64'd5450767261026876886;
    12'd1695: brom_out <= 64'd2359479212055339028;
    12'd1696: brom_out <= 64'd4836003352449041316;
    12'd1697: brom_out <= 64'd6215685832894845107;
    12'd1698: brom_out <= 64'd956565536080223686;
    12'd1699: brom_out <= 64'd3709366288716809584;
    12'd1700: brom_out <= 64'd8051296741047110195;
    12'd1701: brom_out <= 64'd5082200249721761243;
    12'd1702: brom_out <= 64'd4077815017758764724;
    12'd1703: brom_out <= 64'd2646830679214791143;
    12'd1704: brom_out <= 64'd2923414615723271043;
    12'd1705: brom_out <= 64'd9019792797984103029;
    12'd1706: brom_out <= 64'd820027634638271577;
    12'd1707: brom_out <= 64'd2558689606074079344;
    12'd1708: brom_out <= 64'd8026629062288902533;
    12'd1709: brom_out <= 64'd3901615430265803360;
    12'd1710: brom_out <= 64'd2595667101902401433;
    12'd1711: brom_out <= 64'd3645042965713073379;
    12'd1712: brom_out <= 64'd6436331060924184539;
    12'd1713: brom_out <= 64'd5171475373150897937;
    12'd1714: brom_out <= 64'd5549270204663924183;
    12'd1715: brom_out <= 64'd8414575406705992960;
    12'd1716: brom_out <= 64'd6733707155866364304;
    12'd1717: brom_out <= 64'd3582037561619632849;
    12'd1718: brom_out <= 64'd546478178973529773;
    12'd1719: brom_out <= 64'd5586732638848740465;
    12'd1720: brom_out <= 64'd1641922973023157952;
    12'd1721: brom_out <= 64'd815693730606393862;
    12'd1722: brom_out <= 64'd2003304190459111066;
    12'd1723: brom_out <= 64'd7527660023201710545;
    12'd1724: brom_out <= 64'd4681773058202772675;
    12'd1725: brom_out <= 64'd8593145202619771701;
    12'd1726: brom_out <= 64'd3404093846247594996;
    12'd1727: brom_out <= 64'd3486478549657754942;
    12'd1728: brom_out <= 64'd9185509849420767578;
    12'd1729: brom_out <= 64'd6400216294734455669;
    12'd1730: brom_out <= 64'd6282214430396223665;
    12'd1731: brom_out <= 64'd1319517056341783842;
    12'd1732: brom_out <= 64'd6230952056441481807;
    12'd1733: brom_out <= 64'd5263759361851305005;
    12'd1734: brom_out <= 64'd5651215856363377316;
    12'd1735: brom_out <= 64'd1839077451479082854;
    12'd1736: brom_out <= 64'd1546731779372361302;
    12'd1737: brom_out <= 64'd8234108938174010322;
    12'd1738: brom_out <= 64'd3758573853795653427;
    12'd1739: brom_out <= 64'd122506550756017413;
    12'd1740: brom_out <= 64'd1790792280522562723;
    12'd1741: brom_out <= 64'd6466654536513188581;
    12'd1742: brom_out <= 64'd6760985867545539242;
    12'd1743: brom_out <= 64'd8403500667367406851;
    12'd1744: brom_out <= 64'd7995675456769788758;
    12'd1745: brom_out <= 64'd8029507220670853362;
    12'd1746: brom_out <= 64'd3111218648416961668;
    12'd1747: brom_out <= 64'd2521421605044512323;
    12'd1748: brom_out <= 64'd198235807530720187;
    12'd1749: brom_out <= 64'd5152612501000703728;
    12'd1750: brom_out <= 64'd5168690797098687629;
    12'd1751: brom_out <= 64'd1586036392611317199;
    12'd1752: brom_out <= 64'd4849682055056439114;
    12'd1753: brom_out <= 64'd2640079237071612813;
    12'd1754: brom_out <= 64'd1337980060505609637;
    12'd1755: brom_out <= 64'd4740339309841169896;
    12'd1756: brom_out <= 64'd9160052455972965925;
    12'd1757: brom_out <= 64'd3482685859946588622;
    12'd1758: brom_out <= 64'd6411251051681906994;
    12'd1759: brom_out <= 64'd6279407103230115525;
    12'd1760: brom_out <= 64'd9003279055065478956;
    12'd1761: brom_out <= 64'd4849251867203539042;
    12'd1762: brom_out <= 64'd3820044292411662612;
    12'd1763: brom_out <= 64'd2366126602436718469;
    12'd1764: brom_out <= 64'd5011986474190685475;
    12'd1765: brom_out <= 64'd2489326655436610948;
    12'd1766: brom_out <= 64'd8698260697543325537;
    12'd1767: brom_out <= 64'd846810251056707812;
    12'd1768: brom_out <= 64'd869826359180825983;
    12'd1769: brom_out <= 64'd5508432406675787453;
    12'd1770: brom_out <= 64'd3445970765661623385;
    12'd1771: brom_out <= 64'd4183341191108191639;
    12'd1772: brom_out <= 64'd6630229277550940928;
    12'd1773: brom_out <= 64'd1524367001083692685;
    12'd1774: brom_out <= 64'd1664928300054969876;
    12'd1775: brom_out <= 64'd1153272281477598078;
    12'd1776: brom_out <= 64'd1827606411485443129;
    12'd1777: brom_out <= 64'd1892659099199940448;
    12'd1778: brom_out <= 64'd6181880917497703341;
    12'd1779: brom_out <= 64'd1927462247068273250;
    12'd1780: brom_out <= 64'd6949147395764538964;
    12'd1781: brom_out <= 64'd2434856672595838747;
    12'd1782: brom_out <= 64'd7253780654183843384;
    12'd1783: brom_out <= 64'd4643807501097303714;
    12'd1784: brom_out <= 64'd7672998258368931866;
    12'd1785: brom_out <= 64'd166849455930454591;
    12'd1786: brom_out <= 64'd1950822828069733729;
    12'd1787: brom_out <= 64'd1781769378676842139;
    12'd1788: brom_out <= 64'd7530731249570041776;
    12'd1789: brom_out <= 64'd7783916570026358453;
    12'd1790: brom_out <= 64'd8631772682564570593;
    12'd1791: brom_out <= 64'd7708772373098359625;
    12'd1792: brom_out <= 64'd699101306064864663;
    12'd1793: brom_out <= 64'd62383298268607752;
    12'd1794: brom_out <= 64'd7889711590670918676;
    12'd1795: brom_out <= 64'd7816775377648000771;
    12'd1796: brom_out <= 64'd655123889431899961;
    12'd1797: brom_out <= 64'd6822997364396815932;
    12'd1798: brom_out <= 64'd2126660867906687864;
    12'd1799: brom_out <= 64'd7067652521121856833;
    12'd1800: brom_out <= 64'd8219959792660589692;
    12'd1801: brom_out <= 64'd7741423298594687150;
    12'd1802: brom_out <= 64'd8551637415506572346;
    12'd1803: brom_out <= 64'd501434621617250977;
    12'd1804: brom_out <= 64'd8543830174923091154;
    12'd1805: brom_out <= 64'd7799087759160560895;
    12'd1806: brom_out <= 64'd1435047781493708974;
    12'd1807: brom_out <= 64'd1082513074530133782;
    12'd1808: brom_out <= 64'd5893272571222366297;
    12'd1809: brom_out <= 64'd7679327987615867679;
    12'd1810: brom_out <= 64'd7027244046667068898;
    12'd1811: brom_out <= 64'd8516742478246974777;
    12'd1812: brom_out <= 64'd2015889517693822068;
    12'd1813: brom_out <= 64'd8402249683953484293;
    12'd1814: brom_out <= 64'd4971028798941293784;
    12'd1815: brom_out <= 64'd1565712890855058017;
    12'd1816: brom_out <= 64'd4439925312673350003;
    12'd1817: brom_out <= 64'd5876780189316004252;
    12'd1818: brom_out <= 64'd2408543357995828304;
    12'd1819: brom_out <= 64'd4703808339260184091;
    12'd1820: brom_out <= 64'd4798734633597747276;
    12'd1821: brom_out <= 64'd292996083201336963;
    12'd1822: brom_out <= 64'd6781627562122407399;
    12'd1823: brom_out <= 64'd7678224205154604892;
    12'd1824: brom_out <= 64'd69843017785227084;
    12'd1825: brom_out <= 64'd905080829528335056;
    12'd1826: brom_out <= 64'd4891530948138436991;
    12'd1827: brom_out <= 64'd8024688023385731279;
    12'd1828: brom_out <= 64'd8247980103556855667;
    12'd1829: brom_out <= 64'd7549827515419954059;
    12'd1830: brom_out <= 64'd2840283348677403338;
    12'd1831: brom_out <= 64'd7970310816677404075;
    12'd1832: brom_out <= 64'd8225172405297280263;
    12'd1833: brom_out <= 64'd8398591941514173618;
    12'd1834: brom_out <= 64'd7450817543983322844;
    12'd1835: brom_out <= 64'd1851285243088295653;
    12'd1836: brom_out <= 64'd976868090527140556;
    12'd1837: brom_out <= 64'd7186447650655557536;
    12'd1838: brom_out <= 64'd6363705655307338806;
    12'd1839: brom_out <= 64'd2746303970045943107;
    12'd1840: brom_out <= 64'd7645071031480098655;
    12'd1841: brom_out <= 64'd7838092352335735356;
    12'd1842: brom_out <= 64'd3868531777045828691;
    12'd1843: brom_out <= 64'd2506350271925135261;
    12'd1844: brom_out <= 64'd5140288024937627165;
    12'd1845: brom_out <= 64'd1179528608653538977;
    12'd1846: brom_out <= 64'd4538780524597464161;
    12'd1847: brom_out <= 64'd5098416780702440734;
    12'd1848: brom_out <= 64'd5173422508798334624;
    12'd1849: brom_out <= 64'd7068377762402013418;
    12'd1850: brom_out <= 64'd5708860785940369427;
    12'd1851: brom_out <= 64'd3322253652462601701;
    12'd1852: brom_out <= 64'd2600298912569494844;
    12'd1853: brom_out <= 64'd9000423794924863478;
    12'd1854: brom_out <= 64'd6716916671807146392;
    12'd1855: brom_out <= 64'd3079009539254210979;
    12'd1856: brom_out <= 64'd7923677684682802987;
    12'd1857: brom_out <= 64'd9129940191982502832;
    12'd1858: brom_out <= 64'd3815011943812575350;
    12'd1859: brom_out <= 64'd4390475210111465648;
    12'd1860: brom_out <= 64'd2275953281661646751;
    12'd1861: brom_out <= 64'd6075271958765567578;
    12'd1862: brom_out <= 64'd5745260692505968145;
    12'd1863: brom_out <= 64'd797287633007989097;
    12'd1864: brom_out <= 64'd2139689406997953411;
    12'd1865: brom_out <= 64'd902885216720223210;
    12'd1866: brom_out <= 64'd8748419681862114146;
    12'd1867: brom_out <= 64'd2940843062971874248;
    12'd1868: brom_out <= 64'd3729764982569583119;
    12'd1869: brom_out <= 64'd7477596686818285089;
    12'd1870: brom_out <= 64'd1674345919730951813;
    12'd1871: brom_out <= 64'd1900135137736299752;
    12'd1872: brom_out <= 64'd375356035198548383;
    12'd1873: brom_out <= 64'd5954414081382772179;
    12'd1874: brom_out <= 64'd1373369117410510866;
    12'd1875: brom_out <= 64'd874093145357780858;
    12'd1876: brom_out <= 64'd4961919869715327681;
    12'd1877: brom_out <= 64'd6357006725957045398;
    12'd1878: brom_out <= 64'd9052054262515000354;
    12'd1879: brom_out <= 64'd3119795926878188610;
    12'd1880: brom_out <= 64'd511527761999251354;
    12'd1881: brom_out <= 64'd7741012073827083232;
    12'd1882: brom_out <= 64'd3482983880212475854;
    12'd1883: brom_out <= 64'd4946289342964105799;
    12'd1884: brom_out <= 64'd5412893724914022449;
    12'd1885: brom_out <= 64'd2843344465769147130;
    12'd1886: brom_out <= 64'd5032214272686406166;
    12'd1887: brom_out <= 64'd8674281730199549271;
    12'd1888: brom_out <= 64'd5126845061066175356;
    12'd1889: brom_out <= 64'd3530957463225895281;
    12'd1890: brom_out <= 64'd7984550382453767596;
    12'd1891: brom_out <= 64'd1941565973332653447;
    12'd1892: brom_out <= 64'd6181066534637459237;
    12'd1893: brom_out <= 64'd2522950735989919033;
    12'd1894: brom_out <= 64'd8680510475920407927;
    12'd1895: brom_out <= 64'd4928029787718124417;
    12'd1896: brom_out <= 64'd9162350688835803463;
    12'd1897: brom_out <= 64'd4565848593636494677;
    12'd1898: brom_out <= 64'd1414658525045134853;
    12'd1899: brom_out <= 64'd4814867419846616074;
    12'd1900: brom_out <= 64'd841949363898762459;
    12'd1901: brom_out <= 64'd6710867888635545364;
    12'd1902: brom_out <= 64'd486400348447004409;
    12'd1903: brom_out <= 64'd3831753525239012364;
    12'd1904: brom_out <= 64'd796180145389681740;
    12'd1905: brom_out <= 64'd114955450999687352;
    12'd1906: brom_out <= 64'd8371723383654335520;
    12'd1907: brom_out <= 64'd7618198269109257018;
    12'd1908: brom_out <= 64'd6881112568257936145;
    12'd1909: brom_out <= 64'd8154865951547131798;
    12'd1910: brom_out <= 64'd8219861536954301229;
    12'd1911: brom_out <= 64'd6704025482711792486;
    12'd1912: brom_out <= 64'd4119508171639317112;
    12'd1913: brom_out <= 64'd1328025387181652585;
    12'd1914: brom_out <= 64'd2072885801364544572;
    12'd1915: brom_out <= 64'd7266317117570346595;
    12'd1916: brom_out <= 64'd4523573697502160143;
    12'd1917: brom_out <= 64'd2231951319336376728;
    12'd1918: brom_out <= 64'd9096591304164137574;
    12'd1919: brom_out <= 64'd1320547198527024793;
    12'd1920: brom_out <= 64'd1670791095363685175;
    12'd1921: brom_out <= 64'd3917320098766147730;
    12'd1922: brom_out <= 64'd3613147540994151386;
    12'd1923: brom_out <= 64'd7220428068555961202;
    12'd1924: brom_out <= 64'd6268445540391799960;
    12'd1925: brom_out <= 64'd3748546427553799479;
    12'd1926: brom_out <= 64'd333801395018402419;
    12'd1927: brom_out <= 64'd2078333833292311636;
    12'd1928: brom_out <= 64'd5989914729659460893;
    12'd1929: brom_out <= 64'd2080550169979121770;
    12'd1930: brom_out <= 64'd5421197279853390596;
    12'd1931: brom_out <= 64'd3298163028476833569;
    12'd1932: brom_out <= 64'd8498706274306490892;
    12'd1933: brom_out <= 64'd6578345984344235708;
    12'd1934: brom_out <= 64'd7292703967224865486;
    12'd1935: brom_out <= 64'd2984492509020460139;
    12'd1936: brom_out <= 64'd3280526131456603436;
    12'd1937: brom_out <= 64'd7914039759715212288;
    12'd1938: brom_out <= 64'd291195603844344417;
    12'd1939: brom_out <= 64'd5663777043287975940;
    12'd1940: brom_out <= 64'd881381962624186811;
    12'd1941: brom_out <= 64'd3366966051305126938;
    12'd1942: brom_out <= 64'd2351202851047628420;
    12'd1943: brom_out <= 64'd8380172696664431219;
    12'd1944: brom_out <= 64'd3615127351505505023;
    12'd1945: brom_out <= 64'd7870565381825619063;
    12'd1946: brom_out <= 64'd6062993788722341892;
    12'd1947: brom_out <= 64'd2017703862402965552;
    12'd1948: brom_out <= 64'd6148609810148795929;
    12'd1949: brom_out <= 64'd4681885771850953136;
    12'd1950: brom_out <= 64'd599730283692523374;
    12'd1951: brom_out <= 64'd5088451844637495064;
    12'd1952: brom_out <= 64'd8823464365455855293;
    12'd1953: brom_out <= 64'd6261499129228396190;
    12'd1954: brom_out <= 64'd5749262411298578370;
    12'd1955: brom_out <= 64'd5357778098061340193;
    12'd1956: brom_out <= 64'd5139097896322553033;
    12'd1957: brom_out <= 64'd8213543903831367261;
    12'd1958: brom_out <= 64'd8165494333656525134;
    12'd1959: brom_out <= 64'd7997705093244106770;
    12'd1960: brom_out <= 64'd5003529372930301250;
    12'd1961: brom_out <= 64'd6522691292269812797;
    12'd1962: brom_out <= 64'd6319980041019054251;
    12'd1963: brom_out <= 64'd8879506357919806857;
    12'd1964: brom_out <= 64'd3363566323249637328;
    12'd1965: brom_out <= 64'd7901443076583028786;
    12'd1966: brom_out <= 64'd5252122029312962963;
    12'd1967: brom_out <= 64'd1715018151296686515;
    12'd1968: brom_out <= 64'd8323983203612776937;
    12'd1969: brom_out <= 64'd8416441445159376236;
    12'd1970: brom_out <= 64'd2040235830658135393;
    12'd1971: brom_out <= 64'd8480219384681450441;
    12'd1972: brom_out <= 64'd3740576396473059045;
    12'd1973: brom_out <= 64'd2815234299924242613;
    12'd1974: brom_out <= 64'd3289458284692175700;
    12'd1975: brom_out <= 64'd3737566005788852338;
    12'd1976: brom_out <= 64'd5423351720389833865;
    12'd1977: brom_out <= 64'd6669891205375725926;
    12'd1978: brom_out <= 64'd2497038050456785463;
    12'd1979: brom_out <= 64'd8918266820007170405;
    12'd1980: brom_out <= 64'd5408302969401217960;
    12'd1981: brom_out <= 64'd6023400386987486231;
    12'd1982: brom_out <= 64'd7848005646647114461;
    12'd1983: brom_out <= 64'd315347814386475463;
    12'd1984: brom_out <= 64'd228503451388919711;
    12'd1985: brom_out <= 64'd4564125134977115371;
    12'd1986: brom_out <= 64'd2939264214977633037;
    12'd1987: brom_out <= 64'd6822183555527485407;
    12'd1988: brom_out <= 64'd6913883903315781469;
    12'd1989: brom_out <= 64'd7074412356985759977;
    12'd1990: brom_out <= 64'd3506647722126204218;
    12'd1991: brom_out <= 64'd1094028519425961855;
    12'd1992: brom_out <= 64'd498968785704607628;
    12'd1993: brom_out <= 64'd4782115157531486230;
    12'd1994: brom_out <= 64'd911760100456784026;
    12'd1995: brom_out <= 64'd4676447342981270542;
    12'd1996: brom_out <= 64'd3083280881619226755;
    12'd1997: brom_out <= 64'd6602550468570056359;
    12'd1998: brom_out <= 64'd4628098658155976042;
    12'd1999: brom_out <= 64'd5174059410693853581;
    12'd2000: brom_out <= 64'd7002130558985726630;
    12'd2001: brom_out <= 64'd418379368903778945;
    12'd2002: brom_out <= 64'd2804463966393397031;
    12'd2003: brom_out <= 64'd5116562701081850885;
    12'd2004: brom_out <= 64'd3016980039216328962;
    12'd2005: brom_out <= 64'd2296722953695232321;
    12'd2006: brom_out <= 64'd7857926944957203380;
    12'd2007: brom_out <= 64'd7262846507307089798;
    12'd2008: brom_out <= 64'd7471415495952780188;
    12'd2009: brom_out <= 64'd3884405268572847662;
    12'd2010: brom_out <= 64'd713405409942497823;
    12'd2011: brom_out <= 64'd3186532348549307234;
    12'd2012: brom_out <= 64'd9117660520541870682;
    12'd2013: brom_out <= 64'd7094757395937096739;
    12'd2014: brom_out <= 64'd333363560357025169;
    12'd2015: brom_out <= 64'd8065342724630909459;
    12'd2016: brom_out <= 64'd700730835196570872;
    12'd2017: brom_out <= 64'd4797402059262399444;
    12'd2018: brom_out <= 64'd646297118098278772;
    12'd2019: brom_out <= 64'd4563606578771979378;
    12'd2020: brom_out <= 64'd7087203385146507098;
    12'd2021: brom_out <= 64'd498827655396252432;
    12'd2022: brom_out <= 64'd2133757072145401712;
    12'd2023: brom_out <= 64'd6339147614357192038;
    12'd2024: brom_out <= 64'd8584995141337045279;
    12'd2025: brom_out <= 64'd1920532002935580743;
    12'd2026: brom_out <= 64'd830325714398867404;
    12'd2027: brom_out <= 64'd6122157121651334895;
    12'd2028: brom_out <= 64'd6918964554399920495;
    12'd2029: brom_out <= 64'd2077143712079454508;
    12'd2030: brom_out <= 64'd8758553949588800273;
    12'd2031: brom_out <= 64'd25262004549807233;
    12'd2032: brom_out <= 64'd2113561489472542490;
    12'd2033: brom_out <= 64'd5799824691966670023;
    12'd2034: brom_out <= 64'd4130478540001382116;
    12'd2035: brom_out <= 64'd113075564764729104;
    12'd2036: brom_out <= 64'd3835383961103183096;
    12'd2037: brom_out <= 64'd4625028499213347781;
    12'd2038: brom_out <= 64'd2997007021939187347;
    12'd2039: brom_out <= 64'd8461727611525100825;
    12'd2040: brom_out <= 64'd7269045898348823146;
    12'd2041: brom_out <= 64'd5090034518991737864;
    12'd2042: brom_out <= 64'd3031303078308718036;
    12'd2043: brom_out <= 64'd3542987084829734975;
    12'd2044: brom_out <= 64'd8634110784643349010;
    12'd2045: brom_out <= 64'd3528552613765459030;
    12'd2046: brom_out <= 64'd4803548634770013292;
    12'd2047: brom_out <= 64'd9068072491154627648;
    default: brom_out <= 64'h1;
    endcase
end

generate
    if(DELAY == 1) begin
        assign b = brom_out;
    end
endgenerate

endmodule

